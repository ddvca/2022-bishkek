module tm1638_led_display_keys
(
    input   clk,
    input   rst,
    output  tm_clk,
    output  tm_stb,
    inout   tm_dio
);

endmodule
