magic
tech sky130A
magscale 1 2
timestamp 1658639821
<< viali >>
rect 11713 17153 11747 17187
rect 11897 16949 11931 16983
rect 1409 16541 1443 16575
rect 1593 16405 1627 16439
rect 11713 12257 11747 12291
rect 11805 12189 11839 12223
rect 11345 12053 11379 12087
rect 11989 12053 12023 12087
rect 10977 11849 11011 11883
rect 11897 11849 11931 11883
rect 17969 11849 18003 11883
rect 11805 11781 11839 11815
rect 10425 11713 10459 11747
rect 10793 11713 10827 11747
rect 11529 11713 11563 11747
rect 12633 11713 12667 11747
rect 12817 11713 12851 11747
rect 18153 11713 18187 11747
rect 12014 11645 12048 11679
rect 10793 11509 10827 11543
rect 12173 11509 12207 11543
rect 12817 11509 12851 11543
rect 12725 11237 12759 11271
rect 14289 11101 14323 11135
rect 14565 11101 14599 11135
rect 11437 11033 11471 11067
rect 14105 11033 14139 11067
rect 14473 11033 14507 11067
rect 12909 10761 12943 10795
rect 11796 10693 11830 10727
rect 9597 10625 9631 10659
rect 11529 10557 11563 10591
rect 8309 10421 8343 10455
rect 12909 10217 12943 10251
rect 11529 10013 11563 10047
rect 11796 10013 11830 10047
rect 11713 8041 11747 8075
rect 10425 7837 10459 7871
rect 15577 2397 15611 2431
rect 15761 2261 15795 2295
<< metal1 >>
rect 1104 17434 18860 17456
rect 1104 17382 5398 17434
rect 5450 17382 5462 17434
rect 5514 17382 5526 17434
rect 5578 17382 5590 17434
rect 5642 17382 5654 17434
rect 5706 17382 9846 17434
rect 9898 17382 9910 17434
rect 9962 17382 9974 17434
rect 10026 17382 10038 17434
rect 10090 17382 10102 17434
rect 10154 17382 14294 17434
rect 14346 17382 14358 17434
rect 14410 17382 14422 17434
rect 14474 17382 14486 17434
rect 14538 17382 14550 17434
rect 14602 17382 18860 17434
rect 1104 17360 18860 17382
rect 11606 17144 11612 17196
rect 11664 17184 11670 17196
rect 11701 17187 11759 17193
rect 11701 17184 11713 17187
rect 11664 17156 11713 17184
rect 11664 17144 11670 17156
rect 11701 17153 11713 17156
rect 11747 17153 11759 17187
rect 11701 17147 11759 17153
rect 11514 16940 11520 16992
rect 11572 16980 11578 16992
rect 11885 16983 11943 16989
rect 11885 16980 11897 16983
rect 11572 16952 11897 16980
rect 11572 16940 11578 16952
rect 11885 16949 11897 16952
rect 11931 16949 11943 16983
rect 11885 16943 11943 16949
rect 1104 16890 18860 16912
rect 1104 16838 3174 16890
rect 3226 16838 3238 16890
rect 3290 16838 3302 16890
rect 3354 16838 3366 16890
rect 3418 16838 3430 16890
rect 3482 16838 7622 16890
rect 7674 16838 7686 16890
rect 7738 16838 7750 16890
rect 7802 16838 7814 16890
rect 7866 16838 7878 16890
rect 7930 16838 12070 16890
rect 12122 16838 12134 16890
rect 12186 16838 12198 16890
rect 12250 16838 12262 16890
rect 12314 16838 12326 16890
rect 12378 16838 16518 16890
rect 16570 16838 16582 16890
rect 16634 16838 16646 16890
rect 16698 16838 16710 16890
rect 16762 16838 16774 16890
rect 16826 16838 18860 16890
rect 1104 16816 18860 16838
rect 1394 16572 1400 16584
rect 1355 16544 1400 16572
rect 1394 16532 1400 16544
rect 1452 16532 1458 16584
rect 1581 16439 1639 16445
rect 1581 16405 1593 16439
rect 1627 16436 1639 16439
rect 4062 16436 4068 16448
rect 1627 16408 4068 16436
rect 1627 16405 1639 16408
rect 1581 16399 1639 16405
rect 4062 16396 4068 16408
rect 4120 16396 4126 16448
rect 1104 16346 18860 16368
rect 1104 16294 5398 16346
rect 5450 16294 5462 16346
rect 5514 16294 5526 16346
rect 5578 16294 5590 16346
rect 5642 16294 5654 16346
rect 5706 16294 9846 16346
rect 9898 16294 9910 16346
rect 9962 16294 9974 16346
rect 10026 16294 10038 16346
rect 10090 16294 10102 16346
rect 10154 16294 14294 16346
rect 14346 16294 14358 16346
rect 14410 16294 14422 16346
rect 14474 16294 14486 16346
rect 14538 16294 14550 16346
rect 14602 16294 18860 16346
rect 1104 16272 18860 16294
rect 1104 15802 18860 15824
rect 1104 15750 3174 15802
rect 3226 15750 3238 15802
rect 3290 15750 3302 15802
rect 3354 15750 3366 15802
rect 3418 15750 3430 15802
rect 3482 15750 7622 15802
rect 7674 15750 7686 15802
rect 7738 15750 7750 15802
rect 7802 15750 7814 15802
rect 7866 15750 7878 15802
rect 7930 15750 12070 15802
rect 12122 15750 12134 15802
rect 12186 15750 12198 15802
rect 12250 15750 12262 15802
rect 12314 15750 12326 15802
rect 12378 15750 16518 15802
rect 16570 15750 16582 15802
rect 16634 15750 16646 15802
rect 16698 15750 16710 15802
rect 16762 15750 16774 15802
rect 16826 15750 18860 15802
rect 1104 15728 18860 15750
rect 1104 15258 18860 15280
rect 1104 15206 5398 15258
rect 5450 15206 5462 15258
rect 5514 15206 5526 15258
rect 5578 15206 5590 15258
rect 5642 15206 5654 15258
rect 5706 15206 9846 15258
rect 9898 15206 9910 15258
rect 9962 15206 9974 15258
rect 10026 15206 10038 15258
rect 10090 15206 10102 15258
rect 10154 15206 14294 15258
rect 14346 15206 14358 15258
rect 14410 15206 14422 15258
rect 14474 15206 14486 15258
rect 14538 15206 14550 15258
rect 14602 15206 18860 15258
rect 1104 15184 18860 15206
rect 1104 14714 18860 14736
rect 1104 14662 3174 14714
rect 3226 14662 3238 14714
rect 3290 14662 3302 14714
rect 3354 14662 3366 14714
rect 3418 14662 3430 14714
rect 3482 14662 7622 14714
rect 7674 14662 7686 14714
rect 7738 14662 7750 14714
rect 7802 14662 7814 14714
rect 7866 14662 7878 14714
rect 7930 14662 12070 14714
rect 12122 14662 12134 14714
rect 12186 14662 12198 14714
rect 12250 14662 12262 14714
rect 12314 14662 12326 14714
rect 12378 14662 16518 14714
rect 16570 14662 16582 14714
rect 16634 14662 16646 14714
rect 16698 14662 16710 14714
rect 16762 14662 16774 14714
rect 16826 14662 18860 14714
rect 1104 14640 18860 14662
rect 1104 14170 18860 14192
rect 1104 14118 5398 14170
rect 5450 14118 5462 14170
rect 5514 14118 5526 14170
rect 5578 14118 5590 14170
rect 5642 14118 5654 14170
rect 5706 14118 9846 14170
rect 9898 14118 9910 14170
rect 9962 14118 9974 14170
rect 10026 14118 10038 14170
rect 10090 14118 10102 14170
rect 10154 14118 14294 14170
rect 14346 14118 14358 14170
rect 14410 14118 14422 14170
rect 14474 14118 14486 14170
rect 14538 14118 14550 14170
rect 14602 14118 18860 14170
rect 1104 14096 18860 14118
rect 1104 13626 18860 13648
rect 1104 13574 3174 13626
rect 3226 13574 3238 13626
rect 3290 13574 3302 13626
rect 3354 13574 3366 13626
rect 3418 13574 3430 13626
rect 3482 13574 7622 13626
rect 7674 13574 7686 13626
rect 7738 13574 7750 13626
rect 7802 13574 7814 13626
rect 7866 13574 7878 13626
rect 7930 13574 12070 13626
rect 12122 13574 12134 13626
rect 12186 13574 12198 13626
rect 12250 13574 12262 13626
rect 12314 13574 12326 13626
rect 12378 13574 16518 13626
rect 16570 13574 16582 13626
rect 16634 13574 16646 13626
rect 16698 13574 16710 13626
rect 16762 13574 16774 13626
rect 16826 13574 18860 13626
rect 1104 13552 18860 13574
rect 1104 13082 18860 13104
rect 1104 13030 5398 13082
rect 5450 13030 5462 13082
rect 5514 13030 5526 13082
rect 5578 13030 5590 13082
rect 5642 13030 5654 13082
rect 5706 13030 9846 13082
rect 9898 13030 9910 13082
rect 9962 13030 9974 13082
rect 10026 13030 10038 13082
rect 10090 13030 10102 13082
rect 10154 13030 14294 13082
rect 14346 13030 14358 13082
rect 14410 13030 14422 13082
rect 14474 13030 14486 13082
rect 14538 13030 14550 13082
rect 14602 13030 18860 13082
rect 1104 13008 18860 13030
rect 1104 12538 18860 12560
rect 1104 12486 3174 12538
rect 3226 12486 3238 12538
rect 3290 12486 3302 12538
rect 3354 12486 3366 12538
rect 3418 12486 3430 12538
rect 3482 12486 7622 12538
rect 7674 12486 7686 12538
rect 7738 12486 7750 12538
rect 7802 12486 7814 12538
rect 7866 12486 7878 12538
rect 7930 12486 12070 12538
rect 12122 12486 12134 12538
rect 12186 12486 12198 12538
rect 12250 12486 12262 12538
rect 12314 12486 12326 12538
rect 12378 12486 16518 12538
rect 16570 12486 16582 12538
rect 16634 12486 16646 12538
rect 16698 12486 16710 12538
rect 16762 12486 16774 12538
rect 16826 12486 18860 12538
rect 1104 12464 18860 12486
rect 11701 12291 11759 12297
rect 11701 12257 11713 12291
rect 11747 12288 11759 12291
rect 12434 12288 12440 12300
rect 11747 12260 12440 12288
rect 11747 12257 11759 12260
rect 11701 12251 11759 12257
rect 12434 12248 12440 12260
rect 12492 12248 12498 12300
rect 11793 12223 11851 12229
rect 11793 12189 11805 12223
rect 11839 12220 11851 12223
rect 12802 12220 12808 12232
rect 11839 12192 12808 12220
rect 11839 12189 11851 12192
rect 11793 12183 11851 12189
rect 12802 12180 12808 12192
rect 12860 12180 12866 12232
rect 10962 12044 10968 12096
rect 11020 12084 11026 12096
rect 11333 12087 11391 12093
rect 11333 12084 11345 12087
rect 11020 12056 11345 12084
rect 11020 12044 11026 12056
rect 11333 12053 11345 12056
rect 11379 12053 11391 12087
rect 11333 12047 11391 12053
rect 11790 12044 11796 12096
rect 11848 12084 11854 12096
rect 11977 12087 12035 12093
rect 11977 12084 11989 12087
rect 11848 12056 11989 12084
rect 11848 12044 11854 12056
rect 11977 12053 11989 12056
rect 12023 12053 12035 12087
rect 11977 12047 12035 12053
rect 1104 11994 18860 12016
rect 1104 11942 5398 11994
rect 5450 11942 5462 11994
rect 5514 11942 5526 11994
rect 5578 11942 5590 11994
rect 5642 11942 5654 11994
rect 5706 11942 9846 11994
rect 9898 11942 9910 11994
rect 9962 11942 9974 11994
rect 10026 11942 10038 11994
rect 10090 11942 10102 11994
rect 10154 11942 14294 11994
rect 14346 11942 14358 11994
rect 14410 11942 14422 11994
rect 14474 11942 14486 11994
rect 14538 11942 14550 11994
rect 14602 11942 18860 11994
rect 1104 11920 18860 11942
rect 10962 11880 10968 11892
rect 10923 11852 10968 11880
rect 10962 11840 10968 11852
rect 11020 11840 11026 11892
rect 11885 11883 11943 11889
rect 11885 11849 11897 11883
rect 11931 11880 11943 11883
rect 12434 11880 12440 11892
rect 11931 11852 12440 11880
rect 11931 11849 11943 11852
rect 11885 11843 11943 11849
rect 12434 11840 12440 11852
rect 12492 11880 12498 11892
rect 12894 11880 12900 11892
rect 12492 11852 12900 11880
rect 12492 11840 12498 11852
rect 12894 11840 12900 11852
rect 12952 11840 12958 11892
rect 17957 11883 18015 11889
rect 17957 11849 17969 11883
rect 18003 11849 18015 11883
rect 17957 11843 18015 11849
rect 11793 11815 11851 11821
rect 11793 11812 11805 11815
rect 10428 11784 11805 11812
rect 10428 11753 10456 11784
rect 11793 11781 11805 11784
rect 11839 11812 11851 11815
rect 11839 11784 12848 11812
rect 11839 11781 11851 11784
rect 11793 11775 11851 11781
rect 10413 11747 10471 11753
rect 10413 11713 10425 11747
rect 10459 11713 10471 11747
rect 10413 11707 10471 11713
rect 10781 11747 10839 11753
rect 10781 11713 10793 11747
rect 10827 11744 10839 11747
rect 11514 11744 11520 11756
rect 10827 11716 11520 11744
rect 10827 11713 10839 11716
rect 10781 11707 10839 11713
rect 11514 11704 11520 11716
rect 11572 11744 11578 11756
rect 12820 11753 12848 11784
rect 12621 11747 12679 11753
rect 12621 11744 12633 11747
rect 11572 11716 12633 11744
rect 11572 11704 11578 11716
rect 12621 11713 12633 11716
rect 12667 11713 12679 11747
rect 12621 11707 12679 11713
rect 12805 11747 12863 11753
rect 12805 11713 12817 11747
rect 12851 11744 12863 11747
rect 17972 11744 18000 11843
rect 18138 11744 18144 11756
rect 12851 11716 18000 11744
rect 18099 11716 18144 11744
rect 12851 11713 12863 11716
rect 12805 11707 12863 11713
rect 18138 11704 18144 11716
rect 18196 11704 18202 11756
rect 12002 11679 12060 11685
rect 12002 11676 12014 11679
rect 11992 11645 12014 11676
rect 12048 11645 12060 11679
rect 11992 11639 12060 11645
rect 4062 11500 4068 11552
rect 4120 11540 4126 11552
rect 10781 11543 10839 11549
rect 10781 11540 10793 11543
rect 4120 11512 10793 11540
rect 4120 11500 4126 11512
rect 10781 11509 10793 11512
rect 10827 11540 10839 11543
rect 11992 11540 12020 11639
rect 10827 11512 12020 11540
rect 12161 11543 12219 11549
rect 10827 11509 10839 11512
rect 10781 11503 10839 11509
rect 12161 11509 12173 11543
rect 12207 11540 12219 11543
rect 12710 11540 12716 11552
rect 12207 11512 12716 11540
rect 12207 11509 12219 11512
rect 12161 11503 12219 11509
rect 12710 11500 12716 11512
rect 12768 11500 12774 11552
rect 12802 11500 12808 11552
rect 12860 11540 12866 11552
rect 14550 11540 14556 11552
rect 12860 11512 14556 11540
rect 12860 11500 12866 11512
rect 14550 11500 14556 11512
rect 14608 11500 14614 11552
rect 1104 11450 18860 11472
rect 1104 11398 3174 11450
rect 3226 11398 3238 11450
rect 3290 11398 3302 11450
rect 3354 11398 3366 11450
rect 3418 11398 3430 11450
rect 3482 11398 7622 11450
rect 7674 11398 7686 11450
rect 7738 11398 7750 11450
rect 7802 11398 7814 11450
rect 7866 11398 7878 11450
rect 7930 11398 12070 11450
rect 12122 11398 12134 11450
rect 12186 11398 12198 11450
rect 12250 11398 12262 11450
rect 12314 11398 12326 11450
rect 12378 11398 16518 11450
rect 16570 11398 16582 11450
rect 16634 11398 16646 11450
rect 16698 11398 16710 11450
rect 16762 11398 16774 11450
rect 16826 11398 18860 11450
rect 1104 11376 18860 11398
rect 10870 11228 10876 11280
rect 10928 11268 10934 11280
rect 12713 11271 12771 11277
rect 12713 11268 12725 11271
rect 10928 11240 12725 11268
rect 10928 11228 10934 11240
rect 12713 11237 12725 11240
rect 12759 11237 12771 11271
rect 12713 11231 12771 11237
rect 12710 11092 12716 11144
rect 12768 11132 12774 11144
rect 14277 11135 14335 11141
rect 14277 11132 14289 11135
rect 12768 11104 14289 11132
rect 12768 11092 12774 11104
rect 14277 11101 14289 11104
rect 14323 11101 14335 11135
rect 14550 11132 14556 11144
rect 14511 11104 14556 11132
rect 14277 11095 14335 11101
rect 14550 11092 14556 11104
rect 14608 11092 14614 11144
rect 14 11024 20 11076
rect 72 11064 78 11076
rect 11425 11067 11483 11073
rect 11425 11064 11437 11067
rect 72 11036 11437 11064
rect 72 11024 78 11036
rect 11425 11033 11437 11036
rect 11471 11033 11483 11067
rect 11425 11027 11483 11033
rect 12434 11024 12440 11076
rect 12492 11064 12498 11076
rect 14093 11067 14151 11073
rect 14093 11064 14105 11067
rect 12492 11036 14105 11064
rect 12492 11024 12498 11036
rect 14093 11033 14105 11036
rect 14139 11033 14151 11067
rect 14093 11027 14151 11033
rect 14461 11067 14519 11073
rect 14461 11033 14473 11067
rect 14507 11033 14519 11067
rect 14461 11027 14519 11033
rect 13814 10956 13820 11008
rect 13872 10996 13878 11008
rect 14476 10996 14504 11027
rect 15562 10996 15568 11008
rect 13872 10968 15568 10996
rect 13872 10956 13878 10968
rect 15562 10956 15568 10968
rect 15620 10956 15626 11008
rect 1104 10906 18860 10928
rect 1104 10854 5398 10906
rect 5450 10854 5462 10906
rect 5514 10854 5526 10906
rect 5578 10854 5590 10906
rect 5642 10854 5654 10906
rect 5706 10854 9846 10906
rect 9898 10854 9910 10906
rect 9962 10854 9974 10906
rect 10026 10854 10038 10906
rect 10090 10854 10102 10906
rect 10154 10854 14294 10906
rect 14346 10854 14358 10906
rect 14410 10854 14422 10906
rect 14474 10854 14486 10906
rect 14538 10854 14550 10906
rect 14602 10854 18860 10906
rect 1104 10832 18860 10854
rect 12897 10795 12955 10801
rect 12897 10761 12909 10795
rect 12943 10792 12955 10795
rect 13814 10792 13820 10804
rect 12943 10764 13820 10792
rect 12943 10761 12955 10764
rect 12897 10755 12955 10761
rect 13814 10752 13820 10764
rect 13872 10752 13878 10804
rect 11784 10727 11842 10733
rect 11784 10693 11796 10727
rect 11830 10724 11842 10727
rect 12434 10724 12440 10736
rect 11830 10696 12440 10724
rect 11830 10693 11842 10696
rect 11784 10687 11842 10693
rect 12434 10684 12440 10696
rect 12492 10684 12498 10736
rect 9585 10659 9643 10665
rect 9585 10656 9597 10659
rect 9541 10628 9597 10656
rect 9585 10625 9597 10628
rect 9631 10656 9643 10659
rect 10410 10656 10416 10668
rect 9631 10628 10416 10656
rect 9631 10625 9643 10628
rect 9585 10619 9643 10625
rect 10410 10616 10416 10628
rect 10468 10656 10474 10668
rect 10870 10656 10876 10668
rect 10468 10628 10876 10656
rect 10468 10616 10474 10628
rect 10870 10616 10876 10628
rect 10928 10616 10934 10668
rect 11517 10591 11575 10597
rect 11517 10588 11529 10591
rect 9646 10560 11529 10588
rect 8297 10455 8355 10461
rect 8297 10421 8309 10455
rect 8343 10452 8355 10455
rect 9646 10452 9674 10560
rect 11517 10557 11529 10560
rect 11563 10557 11575 10591
rect 11517 10551 11575 10557
rect 8343 10424 9674 10452
rect 8343 10421 8355 10424
rect 8297 10415 8355 10421
rect 1104 10362 18860 10384
rect 1104 10310 3174 10362
rect 3226 10310 3238 10362
rect 3290 10310 3302 10362
rect 3354 10310 3366 10362
rect 3418 10310 3430 10362
rect 3482 10310 7622 10362
rect 7674 10310 7686 10362
rect 7738 10310 7750 10362
rect 7802 10310 7814 10362
rect 7866 10310 7878 10362
rect 7930 10310 12070 10362
rect 12122 10310 12134 10362
rect 12186 10310 12198 10362
rect 12250 10310 12262 10362
rect 12314 10310 12326 10362
rect 12378 10310 16518 10362
rect 16570 10310 16582 10362
rect 16634 10310 16646 10362
rect 16698 10310 16710 10362
rect 16762 10310 16774 10362
rect 16826 10310 18860 10362
rect 1104 10288 18860 10310
rect 12894 10248 12900 10260
rect 12855 10220 12900 10248
rect 12894 10208 12900 10220
rect 12952 10208 12958 10260
rect 11517 10047 11575 10053
rect 11517 10013 11529 10047
rect 11563 10044 11575 10047
rect 11606 10044 11612 10056
rect 11563 10016 11612 10044
rect 11563 10013 11575 10016
rect 11517 10007 11575 10013
rect 11606 10004 11612 10016
rect 11664 10004 11670 10056
rect 11790 10053 11796 10056
rect 11784 10044 11796 10053
rect 11751 10016 11796 10044
rect 11784 10007 11796 10016
rect 11790 10004 11796 10007
rect 11848 10004 11854 10056
rect 1104 9818 18860 9840
rect 1104 9766 5398 9818
rect 5450 9766 5462 9818
rect 5514 9766 5526 9818
rect 5578 9766 5590 9818
rect 5642 9766 5654 9818
rect 5706 9766 9846 9818
rect 9898 9766 9910 9818
rect 9962 9766 9974 9818
rect 10026 9766 10038 9818
rect 10090 9766 10102 9818
rect 10154 9766 14294 9818
rect 14346 9766 14358 9818
rect 14410 9766 14422 9818
rect 14474 9766 14486 9818
rect 14538 9766 14550 9818
rect 14602 9766 18860 9818
rect 1104 9744 18860 9766
rect 1104 9274 18860 9296
rect 1104 9222 3174 9274
rect 3226 9222 3238 9274
rect 3290 9222 3302 9274
rect 3354 9222 3366 9274
rect 3418 9222 3430 9274
rect 3482 9222 7622 9274
rect 7674 9222 7686 9274
rect 7738 9222 7750 9274
rect 7802 9222 7814 9274
rect 7866 9222 7878 9274
rect 7930 9222 12070 9274
rect 12122 9222 12134 9274
rect 12186 9222 12198 9274
rect 12250 9222 12262 9274
rect 12314 9222 12326 9274
rect 12378 9222 16518 9274
rect 16570 9222 16582 9274
rect 16634 9222 16646 9274
rect 16698 9222 16710 9274
rect 16762 9222 16774 9274
rect 16826 9222 18860 9274
rect 1104 9200 18860 9222
rect 1104 8730 18860 8752
rect 1104 8678 5398 8730
rect 5450 8678 5462 8730
rect 5514 8678 5526 8730
rect 5578 8678 5590 8730
rect 5642 8678 5654 8730
rect 5706 8678 9846 8730
rect 9898 8678 9910 8730
rect 9962 8678 9974 8730
rect 10026 8678 10038 8730
rect 10090 8678 10102 8730
rect 10154 8678 14294 8730
rect 14346 8678 14358 8730
rect 14410 8678 14422 8730
rect 14474 8678 14486 8730
rect 14538 8678 14550 8730
rect 14602 8678 18860 8730
rect 1104 8656 18860 8678
rect 1104 8186 18860 8208
rect 1104 8134 3174 8186
rect 3226 8134 3238 8186
rect 3290 8134 3302 8186
rect 3354 8134 3366 8186
rect 3418 8134 3430 8186
rect 3482 8134 7622 8186
rect 7674 8134 7686 8186
rect 7738 8134 7750 8186
rect 7802 8134 7814 8186
rect 7866 8134 7878 8186
rect 7930 8134 12070 8186
rect 12122 8134 12134 8186
rect 12186 8134 12198 8186
rect 12250 8134 12262 8186
rect 12314 8134 12326 8186
rect 12378 8134 16518 8186
rect 16570 8134 16582 8186
rect 16634 8134 16646 8186
rect 16698 8134 16710 8186
rect 16762 8134 16774 8186
rect 16826 8134 18860 8186
rect 1104 8112 18860 8134
rect 11698 8072 11704 8084
rect 11659 8044 11704 8072
rect 11698 8032 11704 8044
rect 11756 8032 11762 8084
rect 10410 7868 10416 7880
rect 10371 7840 10416 7868
rect 10410 7828 10416 7840
rect 10468 7828 10474 7880
rect 1104 7642 18860 7664
rect 1104 7590 5398 7642
rect 5450 7590 5462 7642
rect 5514 7590 5526 7642
rect 5578 7590 5590 7642
rect 5642 7590 5654 7642
rect 5706 7590 9846 7642
rect 9898 7590 9910 7642
rect 9962 7590 9974 7642
rect 10026 7590 10038 7642
rect 10090 7590 10102 7642
rect 10154 7590 14294 7642
rect 14346 7590 14358 7642
rect 14410 7590 14422 7642
rect 14474 7590 14486 7642
rect 14538 7590 14550 7642
rect 14602 7590 18860 7642
rect 1104 7568 18860 7590
rect 1104 7098 18860 7120
rect 1104 7046 3174 7098
rect 3226 7046 3238 7098
rect 3290 7046 3302 7098
rect 3354 7046 3366 7098
rect 3418 7046 3430 7098
rect 3482 7046 7622 7098
rect 7674 7046 7686 7098
rect 7738 7046 7750 7098
rect 7802 7046 7814 7098
rect 7866 7046 7878 7098
rect 7930 7046 12070 7098
rect 12122 7046 12134 7098
rect 12186 7046 12198 7098
rect 12250 7046 12262 7098
rect 12314 7046 12326 7098
rect 12378 7046 16518 7098
rect 16570 7046 16582 7098
rect 16634 7046 16646 7098
rect 16698 7046 16710 7098
rect 16762 7046 16774 7098
rect 16826 7046 18860 7098
rect 1104 7024 18860 7046
rect 1104 6554 18860 6576
rect 1104 6502 5398 6554
rect 5450 6502 5462 6554
rect 5514 6502 5526 6554
rect 5578 6502 5590 6554
rect 5642 6502 5654 6554
rect 5706 6502 9846 6554
rect 9898 6502 9910 6554
rect 9962 6502 9974 6554
rect 10026 6502 10038 6554
rect 10090 6502 10102 6554
rect 10154 6502 14294 6554
rect 14346 6502 14358 6554
rect 14410 6502 14422 6554
rect 14474 6502 14486 6554
rect 14538 6502 14550 6554
rect 14602 6502 18860 6554
rect 1104 6480 18860 6502
rect 1104 6010 18860 6032
rect 1104 5958 3174 6010
rect 3226 5958 3238 6010
rect 3290 5958 3302 6010
rect 3354 5958 3366 6010
rect 3418 5958 3430 6010
rect 3482 5958 7622 6010
rect 7674 5958 7686 6010
rect 7738 5958 7750 6010
rect 7802 5958 7814 6010
rect 7866 5958 7878 6010
rect 7930 5958 12070 6010
rect 12122 5958 12134 6010
rect 12186 5958 12198 6010
rect 12250 5958 12262 6010
rect 12314 5958 12326 6010
rect 12378 5958 16518 6010
rect 16570 5958 16582 6010
rect 16634 5958 16646 6010
rect 16698 5958 16710 6010
rect 16762 5958 16774 6010
rect 16826 5958 18860 6010
rect 1104 5936 18860 5958
rect 1104 5466 18860 5488
rect 1104 5414 5398 5466
rect 5450 5414 5462 5466
rect 5514 5414 5526 5466
rect 5578 5414 5590 5466
rect 5642 5414 5654 5466
rect 5706 5414 9846 5466
rect 9898 5414 9910 5466
rect 9962 5414 9974 5466
rect 10026 5414 10038 5466
rect 10090 5414 10102 5466
rect 10154 5414 14294 5466
rect 14346 5414 14358 5466
rect 14410 5414 14422 5466
rect 14474 5414 14486 5466
rect 14538 5414 14550 5466
rect 14602 5414 18860 5466
rect 1104 5392 18860 5414
rect 1104 4922 18860 4944
rect 1104 4870 3174 4922
rect 3226 4870 3238 4922
rect 3290 4870 3302 4922
rect 3354 4870 3366 4922
rect 3418 4870 3430 4922
rect 3482 4870 7622 4922
rect 7674 4870 7686 4922
rect 7738 4870 7750 4922
rect 7802 4870 7814 4922
rect 7866 4870 7878 4922
rect 7930 4870 12070 4922
rect 12122 4870 12134 4922
rect 12186 4870 12198 4922
rect 12250 4870 12262 4922
rect 12314 4870 12326 4922
rect 12378 4870 16518 4922
rect 16570 4870 16582 4922
rect 16634 4870 16646 4922
rect 16698 4870 16710 4922
rect 16762 4870 16774 4922
rect 16826 4870 18860 4922
rect 1104 4848 18860 4870
rect 1104 4378 18860 4400
rect 1104 4326 5398 4378
rect 5450 4326 5462 4378
rect 5514 4326 5526 4378
rect 5578 4326 5590 4378
rect 5642 4326 5654 4378
rect 5706 4326 9846 4378
rect 9898 4326 9910 4378
rect 9962 4326 9974 4378
rect 10026 4326 10038 4378
rect 10090 4326 10102 4378
rect 10154 4326 14294 4378
rect 14346 4326 14358 4378
rect 14410 4326 14422 4378
rect 14474 4326 14486 4378
rect 14538 4326 14550 4378
rect 14602 4326 18860 4378
rect 1104 4304 18860 4326
rect 1104 3834 18860 3856
rect 1104 3782 3174 3834
rect 3226 3782 3238 3834
rect 3290 3782 3302 3834
rect 3354 3782 3366 3834
rect 3418 3782 3430 3834
rect 3482 3782 7622 3834
rect 7674 3782 7686 3834
rect 7738 3782 7750 3834
rect 7802 3782 7814 3834
rect 7866 3782 7878 3834
rect 7930 3782 12070 3834
rect 12122 3782 12134 3834
rect 12186 3782 12198 3834
rect 12250 3782 12262 3834
rect 12314 3782 12326 3834
rect 12378 3782 16518 3834
rect 16570 3782 16582 3834
rect 16634 3782 16646 3834
rect 16698 3782 16710 3834
rect 16762 3782 16774 3834
rect 16826 3782 18860 3834
rect 1104 3760 18860 3782
rect 1104 3290 18860 3312
rect 1104 3238 5398 3290
rect 5450 3238 5462 3290
rect 5514 3238 5526 3290
rect 5578 3238 5590 3290
rect 5642 3238 5654 3290
rect 5706 3238 9846 3290
rect 9898 3238 9910 3290
rect 9962 3238 9974 3290
rect 10026 3238 10038 3290
rect 10090 3238 10102 3290
rect 10154 3238 14294 3290
rect 14346 3238 14358 3290
rect 14410 3238 14422 3290
rect 14474 3238 14486 3290
rect 14538 3238 14550 3290
rect 14602 3238 18860 3290
rect 1104 3216 18860 3238
rect 1104 2746 18860 2768
rect 1104 2694 3174 2746
rect 3226 2694 3238 2746
rect 3290 2694 3302 2746
rect 3354 2694 3366 2746
rect 3418 2694 3430 2746
rect 3482 2694 7622 2746
rect 7674 2694 7686 2746
rect 7738 2694 7750 2746
rect 7802 2694 7814 2746
rect 7866 2694 7878 2746
rect 7930 2694 12070 2746
rect 12122 2694 12134 2746
rect 12186 2694 12198 2746
rect 12250 2694 12262 2746
rect 12314 2694 12326 2746
rect 12378 2694 16518 2746
rect 16570 2694 16582 2746
rect 16634 2694 16646 2746
rect 16698 2694 16710 2746
rect 16762 2694 16774 2746
rect 16826 2694 18860 2746
rect 1104 2672 18860 2694
rect 15562 2428 15568 2440
rect 15523 2400 15568 2428
rect 15562 2388 15568 2400
rect 15620 2388 15626 2440
rect 15470 2252 15476 2304
rect 15528 2292 15534 2304
rect 15749 2295 15807 2301
rect 15749 2292 15761 2295
rect 15528 2264 15761 2292
rect 15528 2252 15534 2264
rect 15749 2261 15761 2264
rect 15795 2261 15807 2295
rect 15749 2255 15807 2261
rect 1104 2202 18860 2224
rect 1104 2150 5398 2202
rect 5450 2150 5462 2202
rect 5514 2150 5526 2202
rect 5578 2150 5590 2202
rect 5642 2150 5654 2202
rect 5706 2150 9846 2202
rect 9898 2150 9910 2202
rect 9962 2150 9974 2202
rect 10026 2150 10038 2202
rect 10090 2150 10102 2202
rect 10154 2150 14294 2202
rect 14346 2150 14358 2202
rect 14410 2150 14422 2202
rect 14474 2150 14486 2202
rect 14538 2150 14550 2202
rect 14602 2150 18860 2202
rect 1104 2128 18860 2150
<< via1 >>
rect 5398 17382 5450 17434
rect 5462 17382 5514 17434
rect 5526 17382 5578 17434
rect 5590 17382 5642 17434
rect 5654 17382 5706 17434
rect 9846 17382 9898 17434
rect 9910 17382 9962 17434
rect 9974 17382 10026 17434
rect 10038 17382 10090 17434
rect 10102 17382 10154 17434
rect 14294 17382 14346 17434
rect 14358 17382 14410 17434
rect 14422 17382 14474 17434
rect 14486 17382 14538 17434
rect 14550 17382 14602 17434
rect 11612 17144 11664 17196
rect 11520 16940 11572 16992
rect 3174 16838 3226 16890
rect 3238 16838 3290 16890
rect 3302 16838 3354 16890
rect 3366 16838 3418 16890
rect 3430 16838 3482 16890
rect 7622 16838 7674 16890
rect 7686 16838 7738 16890
rect 7750 16838 7802 16890
rect 7814 16838 7866 16890
rect 7878 16838 7930 16890
rect 12070 16838 12122 16890
rect 12134 16838 12186 16890
rect 12198 16838 12250 16890
rect 12262 16838 12314 16890
rect 12326 16838 12378 16890
rect 16518 16838 16570 16890
rect 16582 16838 16634 16890
rect 16646 16838 16698 16890
rect 16710 16838 16762 16890
rect 16774 16838 16826 16890
rect 1400 16575 1452 16584
rect 1400 16541 1409 16575
rect 1409 16541 1443 16575
rect 1443 16541 1452 16575
rect 1400 16532 1452 16541
rect 4068 16396 4120 16448
rect 5398 16294 5450 16346
rect 5462 16294 5514 16346
rect 5526 16294 5578 16346
rect 5590 16294 5642 16346
rect 5654 16294 5706 16346
rect 9846 16294 9898 16346
rect 9910 16294 9962 16346
rect 9974 16294 10026 16346
rect 10038 16294 10090 16346
rect 10102 16294 10154 16346
rect 14294 16294 14346 16346
rect 14358 16294 14410 16346
rect 14422 16294 14474 16346
rect 14486 16294 14538 16346
rect 14550 16294 14602 16346
rect 3174 15750 3226 15802
rect 3238 15750 3290 15802
rect 3302 15750 3354 15802
rect 3366 15750 3418 15802
rect 3430 15750 3482 15802
rect 7622 15750 7674 15802
rect 7686 15750 7738 15802
rect 7750 15750 7802 15802
rect 7814 15750 7866 15802
rect 7878 15750 7930 15802
rect 12070 15750 12122 15802
rect 12134 15750 12186 15802
rect 12198 15750 12250 15802
rect 12262 15750 12314 15802
rect 12326 15750 12378 15802
rect 16518 15750 16570 15802
rect 16582 15750 16634 15802
rect 16646 15750 16698 15802
rect 16710 15750 16762 15802
rect 16774 15750 16826 15802
rect 5398 15206 5450 15258
rect 5462 15206 5514 15258
rect 5526 15206 5578 15258
rect 5590 15206 5642 15258
rect 5654 15206 5706 15258
rect 9846 15206 9898 15258
rect 9910 15206 9962 15258
rect 9974 15206 10026 15258
rect 10038 15206 10090 15258
rect 10102 15206 10154 15258
rect 14294 15206 14346 15258
rect 14358 15206 14410 15258
rect 14422 15206 14474 15258
rect 14486 15206 14538 15258
rect 14550 15206 14602 15258
rect 3174 14662 3226 14714
rect 3238 14662 3290 14714
rect 3302 14662 3354 14714
rect 3366 14662 3418 14714
rect 3430 14662 3482 14714
rect 7622 14662 7674 14714
rect 7686 14662 7738 14714
rect 7750 14662 7802 14714
rect 7814 14662 7866 14714
rect 7878 14662 7930 14714
rect 12070 14662 12122 14714
rect 12134 14662 12186 14714
rect 12198 14662 12250 14714
rect 12262 14662 12314 14714
rect 12326 14662 12378 14714
rect 16518 14662 16570 14714
rect 16582 14662 16634 14714
rect 16646 14662 16698 14714
rect 16710 14662 16762 14714
rect 16774 14662 16826 14714
rect 5398 14118 5450 14170
rect 5462 14118 5514 14170
rect 5526 14118 5578 14170
rect 5590 14118 5642 14170
rect 5654 14118 5706 14170
rect 9846 14118 9898 14170
rect 9910 14118 9962 14170
rect 9974 14118 10026 14170
rect 10038 14118 10090 14170
rect 10102 14118 10154 14170
rect 14294 14118 14346 14170
rect 14358 14118 14410 14170
rect 14422 14118 14474 14170
rect 14486 14118 14538 14170
rect 14550 14118 14602 14170
rect 3174 13574 3226 13626
rect 3238 13574 3290 13626
rect 3302 13574 3354 13626
rect 3366 13574 3418 13626
rect 3430 13574 3482 13626
rect 7622 13574 7674 13626
rect 7686 13574 7738 13626
rect 7750 13574 7802 13626
rect 7814 13574 7866 13626
rect 7878 13574 7930 13626
rect 12070 13574 12122 13626
rect 12134 13574 12186 13626
rect 12198 13574 12250 13626
rect 12262 13574 12314 13626
rect 12326 13574 12378 13626
rect 16518 13574 16570 13626
rect 16582 13574 16634 13626
rect 16646 13574 16698 13626
rect 16710 13574 16762 13626
rect 16774 13574 16826 13626
rect 5398 13030 5450 13082
rect 5462 13030 5514 13082
rect 5526 13030 5578 13082
rect 5590 13030 5642 13082
rect 5654 13030 5706 13082
rect 9846 13030 9898 13082
rect 9910 13030 9962 13082
rect 9974 13030 10026 13082
rect 10038 13030 10090 13082
rect 10102 13030 10154 13082
rect 14294 13030 14346 13082
rect 14358 13030 14410 13082
rect 14422 13030 14474 13082
rect 14486 13030 14538 13082
rect 14550 13030 14602 13082
rect 3174 12486 3226 12538
rect 3238 12486 3290 12538
rect 3302 12486 3354 12538
rect 3366 12486 3418 12538
rect 3430 12486 3482 12538
rect 7622 12486 7674 12538
rect 7686 12486 7738 12538
rect 7750 12486 7802 12538
rect 7814 12486 7866 12538
rect 7878 12486 7930 12538
rect 12070 12486 12122 12538
rect 12134 12486 12186 12538
rect 12198 12486 12250 12538
rect 12262 12486 12314 12538
rect 12326 12486 12378 12538
rect 16518 12486 16570 12538
rect 16582 12486 16634 12538
rect 16646 12486 16698 12538
rect 16710 12486 16762 12538
rect 16774 12486 16826 12538
rect 12440 12248 12492 12300
rect 12808 12180 12860 12232
rect 10968 12044 11020 12096
rect 11796 12044 11848 12096
rect 5398 11942 5450 11994
rect 5462 11942 5514 11994
rect 5526 11942 5578 11994
rect 5590 11942 5642 11994
rect 5654 11942 5706 11994
rect 9846 11942 9898 11994
rect 9910 11942 9962 11994
rect 9974 11942 10026 11994
rect 10038 11942 10090 11994
rect 10102 11942 10154 11994
rect 14294 11942 14346 11994
rect 14358 11942 14410 11994
rect 14422 11942 14474 11994
rect 14486 11942 14538 11994
rect 14550 11942 14602 11994
rect 10968 11883 11020 11892
rect 10968 11849 10977 11883
rect 10977 11849 11011 11883
rect 11011 11849 11020 11883
rect 10968 11840 11020 11849
rect 12440 11840 12492 11892
rect 12900 11840 12952 11892
rect 11520 11747 11572 11756
rect 11520 11713 11529 11747
rect 11529 11713 11563 11747
rect 11563 11713 11572 11747
rect 11520 11704 11572 11713
rect 18144 11747 18196 11756
rect 18144 11713 18153 11747
rect 18153 11713 18187 11747
rect 18187 11713 18196 11747
rect 18144 11704 18196 11713
rect 4068 11500 4120 11552
rect 12716 11500 12768 11552
rect 12808 11543 12860 11552
rect 12808 11509 12817 11543
rect 12817 11509 12851 11543
rect 12851 11509 12860 11543
rect 12808 11500 12860 11509
rect 14556 11500 14608 11552
rect 3174 11398 3226 11450
rect 3238 11398 3290 11450
rect 3302 11398 3354 11450
rect 3366 11398 3418 11450
rect 3430 11398 3482 11450
rect 7622 11398 7674 11450
rect 7686 11398 7738 11450
rect 7750 11398 7802 11450
rect 7814 11398 7866 11450
rect 7878 11398 7930 11450
rect 12070 11398 12122 11450
rect 12134 11398 12186 11450
rect 12198 11398 12250 11450
rect 12262 11398 12314 11450
rect 12326 11398 12378 11450
rect 16518 11398 16570 11450
rect 16582 11398 16634 11450
rect 16646 11398 16698 11450
rect 16710 11398 16762 11450
rect 16774 11398 16826 11450
rect 10876 11228 10928 11280
rect 12716 11092 12768 11144
rect 14556 11135 14608 11144
rect 14556 11101 14565 11135
rect 14565 11101 14599 11135
rect 14599 11101 14608 11135
rect 14556 11092 14608 11101
rect 20 11024 72 11076
rect 12440 11024 12492 11076
rect 13820 10956 13872 11008
rect 15568 10956 15620 11008
rect 5398 10854 5450 10906
rect 5462 10854 5514 10906
rect 5526 10854 5578 10906
rect 5590 10854 5642 10906
rect 5654 10854 5706 10906
rect 9846 10854 9898 10906
rect 9910 10854 9962 10906
rect 9974 10854 10026 10906
rect 10038 10854 10090 10906
rect 10102 10854 10154 10906
rect 14294 10854 14346 10906
rect 14358 10854 14410 10906
rect 14422 10854 14474 10906
rect 14486 10854 14538 10906
rect 14550 10854 14602 10906
rect 13820 10752 13872 10804
rect 12440 10684 12492 10736
rect 10416 10616 10468 10668
rect 10876 10616 10928 10668
rect 3174 10310 3226 10362
rect 3238 10310 3290 10362
rect 3302 10310 3354 10362
rect 3366 10310 3418 10362
rect 3430 10310 3482 10362
rect 7622 10310 7674 10362
rect 7686 10310 7738 10362
rect 7750 10310 7802 10362
rect 7814 10310 7866 10362
rect 7878 10310 7930 10362
rect 12070 10310 12122 10362
rect 12134 10310 12186 10362
rect 12198 10310 12250 10362
rect 12262 10310 12314 10362
rect 12326 10310 12378 10362
rect 16518 10310 16570 10362
rect 16582 10310 16634 10362
rect 16646 10310 16698 10362
rect 16710 10310 16762 10362
rect 16774 10310 16826 10362
rect 12900 10251 12952 10260
rect 12900 10217 12909 10251
rect 12909 10217 12943 10251
rect 12943 10217 12952 10251
rect 12900 10208 12952 10217
rect 11612 10004 11664 10056
rect 11796 10047 11848 10056
rect 11796 10013 11830 10047
rect 11830 10013 11848 10047
rect 11796 10004 11848 10013
rect 5398 9766 5450 9818
rect 5462 9766 5514 9818
rect 5526 9766 5578 9818
rect 5590 9766 5642 9818
rect 5654 9766 5706 9818
rect 9846 9766 9898 9818
rect 9910 9766 9962 9818
rect 9974 9766 10026 9818
rect 10038 9766 10090 9818
rect 10102 9766 10154 9818
rect 14294 9766 14346 9818
rect 14358 9766 14410 9818
rect 14422 9766 14474 9818
rect 14486 9766 14538 9818
rect 14550 9766 14602 9818
rect 3174 9222 3226 9274
rect 3238 9222 3290 9274
rect 3302 9222 3354 9274
rect 3366 9222 3418 9274
rect 3430 9222 3482 9274
rect 7622 9222 7674 9274
rect 7686 9222 7738 9274
rect 7750 9222 7802 9274
rect 7814 9222 7866 9274
rect 7878 9222 7930 9274
rect 12070 9222 12122 9274
rect 12134 9222 12186 9274
rect 12198 9222 12250 9274
rect 12262 9222 12314 9274
rect 12326 9222 12378 9274
rect 16518 9222 16570 9274
rect 16582 9222 16634 9274
rect 16646 9222 16698 9274
rect 16710 9222 16762 9274
rect 16774 9222 16826 9274
rect 5398 8678 5450 8730
rect 5462 8678 5514 8730
rect 5526 8678 5578 8730
rect 5590 8678 5642 8730
rect 5654 8678 5706 8730
rect 9846 8678 9898 8730
rect 9910 8678 9962 8730
rect 9974 8678 10026 8730
rect 10038 8678 10090 8730
rect 10102 8678 10154 8730
rect 14294 8678 14346 8730
rect 14358 8678 14410 8730
rect 14422 8678 14474 8730
rect 14486 8678 14538 8730
rect 14550 8678 14602 8730
rect 3174 8134 3226 8186
rect 3238 8134 3290 8186
rect 3302 8134 3354 8186
rect 3366 8134 3418 8186
rect 3430 8134 3482 8186
rect 7622 8134 7674 8186
rect 7686 8134 7738 8186
rect 7750 8134 7802 8186
rect 7814 8134 7866 8186
rect 7878 8134 7930 8186
rect 12070 8134 12122 8186
rect 12134 8134 12186 8186
rect 12198 8134 12250 8186
rect 12262 8134 12314 8186
rect 12326 8134 12378 8186
rect 16518 8134 16570 8186
rect 16582 8134 16634 8186
rect 16646 8134 16698 8186
rect 16710 8134 16762 8186
rect 16774 8134 16826 8186
rect 11704 8075 11756 8084
rect 11704 8041 11713 8075
rect 11713 8041 11747 8075
rect 11747 8041 11756 8075
rect 11704 8032 11756 8041
rect 10416 7871 10468 7880
rect 10416 7837 10425 7871
rect 10425 7837 10459 7871
rect 10459 7837 10468 7871
rect 10416 7828 10468 7837
rect 5398 7590 5450 7642
rect 5462 7590 5514 7642
rect 5526 7590 5578 7642
rect 5590 7590 5642 7642
rect 5654 7590 5706 7642
rect 9846 7590 9898 7642
rect 9910 7590 9962 7642
rect 9974 7590 10026 7642
rect 10038 7590 10090 7642
rect 10102 7590 10154 7642
rect 14294 7590 14346 7642
rect 14358 7590 14410 7642
rect 14422 7590 14474 7642
rect 14486 7590 14538 7642
rect 14550 7590 14602 7642
rect 3174 7046 3226 7098
rect 3238 7046 3290 7098
rect 3302 7046 3354 7098
rect 3366 7046 3418 7098
rect 3430 7046 3482 7098
rect 7622 7046 7674 7098
rect 7686 7046 7738 7098
rect 7750 7046 7802 7098
rect 7814 7046 7866 7098
rect 7878 7046 7930 7098
rect 12070 7046 12122 7098
rect 12134 7046 12186 7098
rect 12198 7046 12250 7098
rect 12262 7046 12314 7098
rect 12326 7046 12378 7098
rect 16518 7046 16570 7098
rect 16582 7046 16634 7098
rect 16646 7046 16698 7098
rect 16710 7046 16762 7098
rect 16774 7046 16826 7098
rect 5398 6502 5450 6554
rect 5462 6502 5514 6554
rect 5526 6502 5578 6554
rect 5590 6502 5642 6554
rect 5654 6502 5706 6554
rect 9846 6502 9898 6554
rect 9910 6502 9962 6554
rect 9974 6502 10026 6554
rect 10038 6502 10090 6554
rect 10102 6502 10154 6554
rect 14294 6502 14346 6554
rect 14358 6502 14410 6554
rect 14422 6502 14474 6554
rect 14486 6502 14538 6554
rect 14550 6502 14602 6554
rect 3174 5958 3226 6010
rect 3238 5958 3290 6010
rect 3302 5958 3354 6010
rect 3366 5958 3418 6010
rect 3430 5958 3482 6010
rect 7622 5958 7674 6010
rect 7686 5958 7738 6010
rect 7750 5958 7802 6010
rect 7814 5958 7866 6010
rect 7878 5958 7930 6010
rect 12070 5958 12122 6010
rect 12134 5958 12186 6010
rect 12198 5958 12250 6010
rect 12262 5958 12314 6010
rect 12326 5958 12378 6010
rect 16518 5958 16570 6010
rect 16582 5958 16634 6010
rect 16646 5958 16698 6010
rect 16710 5958 16762 6010
rect 16774 5958 16826 6010
rect 5398 5414 5450 5466
rect 5462 5414 5514 5466
rect 5526 5414 5578 5466
rect 5590 5414 5642 5466
rect 5654 5414 5706 5466
rect 9846 5414 9898 5466
rect 9910 5414 9962 5466
rect 9974 5414 10026 5466
rect 10038 5414 10090 5466
rect 10102 5414 10154 5466
rect 14294 5414 14346 5466
rect 14358 5414 14410 5466
rect 14422 5414 14474 5466
rect 14486 5414 14538 5466
rect 14550 5414 14602 5466
rect 3174 4870 3226 4922
rect 3238 4870 3290 4922
rect 3302 4870 3354 4922
rect 3366 4870 3418 4922
rect 3430 4870 3482 4922
rect 7622 4870 7674 4922
rect 7686 4870 7738 4922
rect 7750 4870 7802 4922
rect 7814 4870 7866 4922
rect 7878 4870 7930 4922
rect 12070 4870 12122 4922
rect 12134 4870 12186 4922
rect 12198 4870 12250 4922
rect 12262 4870 12314 4922
rect 12326 4870 12378 4922
rect 16518 4870 16570 4922
rect 16582 4870 16634 4922
rect 16646 4870 16698 4922
rect 16710 4870 16762 4922
rect 16774 4870 16826 4922
rect 5398 4326 5450 4378
rect 5462 4326 5514 4378
rect 5526 4326 5578 4378
rect 5590 4326 5642 4378
rect 5654 4326 5706 4378
rect 9846 4326 9898 4378
rect 9910 4326 9962 4378
rect 9974 4326 10026 4378
rect 10038 4326 10090 4378
rect 10102 4326 10154 4378
rect 14294 4326 14346 4378
rect 14358 4326 14410 4378
rect 14422 4326 14474 4378
rect 14486 4326 14538 4378
rect 14550 4326 14602 4378
rect 3174 3782 3226 3834
rect 3238 3782 3290 3834
rect 3302 3782 3354 3834
rect 3366 3782 3418 3834
rect 3430 3782 3482 3834
rect 7622 3782 7674 3834
rect 7686 3782 7738 3834
rect 7750 3782 7802 3834
rect 7814 3782 7866 3834
rect 7878 3782 7930 3834
rect 12070 3782 12122 3834
rect 12134 3782 12186 3834
rect 12198 3782 12250 3834
rect 12262 3782 12314 3834
rect 12326 3782 12378 3834
rect 16518 3782 16570 3834
rect 16582 3782 16634 3834
rect 16646 3782 16698 3834
rect 16710 3782 16762 3834
rect 16774 3782 16826 3834
rect 5398 3238 5450 3290
rect 5462 3238 5514 3290
rect 5526 3238 5578 3290
rect 5590 3238 5642 3290
rect 5654 3238 5706 3290
rect 9846 3238 9898 3290
rect 9910 3238 9962 3290
rect 9974 3238 10026 3290
rect 10038 3238 10090 3290
rect 10102 3238 10154 3290
rect 14294 3238 14346 3290
rect 14358 3238 14410 3290
rect 14422 3238 14474 3290
rect 14486 3238 14538 3290
rect 14550 3238 14602 3290
rect 3174 2694 3226 2746
rect 3238 2694 3290 2746
rect 3302 2694 3354 2746
rect 3366 2694 3418 2746
rect 3430 2694 3482 2746
rect 7622 2694 7674 2746
rect 7686 2694 7738 2746
rect 7750 2694 7802 2746
rect 7814 2694 7866 2746
rect 7878 2694 7930 2746
rect 12070 2694 12122 2746
rect 12134 2694 12186 2746
rect 12198 2694 12250 2746
rect 12262 2694 12314 2746
rect 12326 2694 12378 2746
rect 16518 2694 16570 2746
rect 16582 2694 16634 2746
rect 16646 2694 16698 2746
rect 16710 2694 16762 2746
rect 16774 2694 16826 2746
rect 15568 2431 15620 2440
rect 15568 2397 15577 2431
rect 15577 2397 15611 2431
rect 15611 2397 15620 2431
rect 15568 2388 15620 2397
rect 15476 2252 15528 2304
rect 5398 2150 5450 2202
rect 5462 2150 5514 2202
rect 5526 2150 5578 2202
rect 5590 2150 5642 2202
rect 5654 2150 5706 2202
rect 9846 2150 9898 2202
rect 9910 2150 9962 2202
rect 9974 2150 10026 2202
rect 10038 2150 10090 2202
rect 10102 2150 10154 2202
rect 14294 2150 14346 2202
rect 14358 2150 14410 2202
rect 14422 2150 14474 2202
rect 14486 2150 14538 2202
rect 14550 2150 14602 2202
<< metal2 >>
rect 11610 19200 11666 20000
rect 5398 17436 5706 17445
rect 5398 17434 5404 17436
rect 5460 17434 5484 17436
rect 5540 17434 5564 17436
rect 5620 17434 5644 17436
rect 5700 17434 5706 17436
rect 5460 17382 5462 17434
rect 5642 17382 5644 17434
rect 5398 17380 5404 17382
rect 5460 17380 5484 17382
rect 5540 17380 5564 17382
rect 5620 17380 5644 17382
rect 5700 17380 5706 17382
rect 5398 17371 5706 17380
rect 9846 17436 10154 17445
rect 9846 17434 9852 17436
rect 9908 17434 9932 17436
rect 9988 17434 10012 17436
rect 10068 17434 10092 17436
rect 10148 17434 10154 17436
rect 9908 17382 9910 17434
rect 10090 17382 10092 17434
rect 9846 17380 9852 17382
rect 9908 17380 9932 17382
rect 9988 17380 10012 17382
rect 10068 17380 10092 17382
rect 10148 17380 10154 17382
rect 9846 17371 10154 17380
rect 11624 17202 11652 19200
rect 14294 17436 14602 17445
rect 14294 17434 14300 17436
rect 14356 17434 14380 17436
rect 14436 17434 14460 17436
rect 14516 17434 14540 17436
rect 14596 17434 14602 17436
rect 14356 17382 14358 17434
rect 14538 17382 14540 17434
rect 14294 17380 14300 17382
rect 14356 17380 14380 17382
rect 14436 17380 14460 17382
rect 14516 17380 14540 17382
rect 14596 17380 14602 17382
rect 14294 17371 14602 17380
rect 11612 17196 11664 17202
rect 11612 17138 11664 17144
rect 11520 16992 11572 16998
rect 11520 16934 11572 16940
rect 3174 16892 3482 16901
rect 3174 16890 3180 16892
rect 3236 16890 3260 16892
rect 3316 16890 3340 16892
rect 3396 16890 3420 16892
rect 3476 16890 3482 16892
rect 3236 16838 3238 16890
rect 3418 16838 3420 16890
rect 3174 16836 3180 16838
rect 3236 16836 3260 16838
rect 3316 16836 3340 16838
rect 3396 16836 3420 16838
rect 3476 16836 3482 16838
rect 3174 16827 3482 16836
rect 7622 16892 7930 16901
rect 7622 16890 7628 16892
rect 7684 16890 7708 16892
rect 7764 16890 7788 16892
rect 7844 16890 7868 16892
rect 7924 16890 7930 16892
rect 7684 16838 7686 16890
rect 7866 16838 7868 16890
rect 7622 16836 7628 16838
rect 7684 16836 7708 16838
rect 7764 16836 7788 16838
rect 7844 16836 7868 16838
rect 7924 16836 7930 16838
rect 7622 16827 7930 16836
rect 1400 16584 1452 16590
rect 1400 16526 1452 16532
rect 1412 16425 1440 16526
rect 4068 16448 4120 16454
rect 1398 16416 1454 16425
rect 4068 16390 4120 16396
rect 1398 16351 1454 16360
rect 3174 15804 3482 15813
rect 3174 15802 3180 15804
rect 3236 15802 3260 15804
rect 3316 15802 3340 15804
rect 3396 15802 3420 15804
rect 3476 15802 3482 15804
rect 3236 15750 3238 15802
rect 3418 15750 3420 15802
rect 3174 15748 3180 15750
rect 3236 15748 3260 15750
rect 3316 15748 3340 15750
rect 3396 15748 3420 15750
rect 3476 15748 3482 15750
rect 3174 15739 3482 15748
rect 3174 14716 3482 14725
rect 3174 14714 3180 14716
rect 3236 14714 3260 14716
rect 3316 14714 3340 14716
rect 3396 14714 3420 14716
rect 3476 14714 3482 14716
rect 3236 14662 3238 14714
rect 3418 14662 3420 14714
rect 3174 14660 3180 14662
rect 3236 14660 3260 14662
rect 3316 14660 3340 14662
rect 3396 14660 3420 14662
rect 3476 14660 3482 14662
rect 3174 14651 3482 14660
rect 3174 13628 3482 13637
rect 3174 13626 3180 13628
rect 3236 13626 3260 13628
rect 3316 13626 3340 13628
rect 3396 13626 3420 13628
rect 3476 13626 3482 13628
rect 3236 13574 3238 13626
rect 3418 13574 3420 13626
rect 3174 13572 3180 13574
rect 3236 13572 3260 13574
rect 3316 13572 3340 13574
rect 3396 13572 3420 13574
rect 3476 13572 3482 13574
rect 3174 13563 3482 13572
rect 3174 12540 3482 12549
rect 3174 12538 3180 12540
rect 3236 12538 3260 12540
rect 3316 12538 3340 12540
rect 3396 12538 3420 12540
rect 3476 12538 3482 12540
rect 3236 12486 3238 12538
rect 3418 12486 3420 12538
rect 3174 12484 3180 12486
rect 3236 12484 3260 12486
rect 3316 12484 3340 12486
rect 3396 12484 3420 12486
rect 3476 12484 3482 12486
rect 3174 12475 3482 12484
rect 4080 11558 4108 16390
rect 5398 16348 5706 16357
rect 5398 16346 5404 16348
rect 5460 16346 5484 16348
rect 5540 16346 5564 16348
rect 5620 16346 5644 16348
rect 5700 16346 5706 16348
rect 5460 16294 5462 16346
rect 5642 16294 5644 16346
rect 5398 16292 5404 16294
rect 5460 16292 5484 16294
rect 5540 16292 5564 16294
rect 5620 16292 5644 16294
rect 5700 16292 5706 16294
rect 5398 16283 5706 16292
rect 9846 16348 10154 16357
rect 9846 16346 9852 16348
rect 9908 16346 9932 16348
rect 9988 16346 10012 16348
rect 10068 16346 10092 16348
rect 10148 16346 10154 16348
rect 9908 16294 9910 16346
rect 10090 16294 10092 16346
rect 9846 16292 9852 16294
rect 9908 16292 9932 16294
rect 9988 16292 10012 16294
rect 10068 16292 10092 16294
rect 10148 16292 10154 16294
rect 9846 16283 10154 16292
rect 7622 15804 7930 15813
rect 7622 15802 7628 15804
rect 7684 15802 7708 15804
rect 7764 15802 7788 15804
rect 7844 15802 7868 15804
rect 7924 15802 7930 15804
rect 7684 15750 7686 15802
rect 7866 15750 7868 15802
rect 7622 15748 7628 15750
rect 7684 15748 7708 15750
rect 7764 15748 7788 15750
rect 7844 15748 7868 15750
rect 7924 15748 7930 15750
rect 7622 15739 7930 15748
rect 5398 15260 5706 15269
rect 5398 15258 5404 15260
rect 5460 15258 5484 15260
rect 5540 15258 5564 15260
rect 5620 15258 5644 15260
rect 5700 15258 5706 15260
rect 5460 15206 5462 15258
rect 5642 15206 5644 15258
rect 5398 15204 5404 15206
rect 5460 15204 5484 15206
rect 5540 15204 5564 15206
rect 5620 15204 5644 15206
rect 5700 15204 5706 15206
rect 5398 15195 5706 15204
rect 9846 15260 10154 15269
rect 9846 15258 9852 15260
rect 9908 15258 9932 15260
rect 9988 15258 10012 15260
rect 10068 15258 10092 15260
rect 10148 15258 10154 15260
rect 9908 15206 9910 15258
rect 10090 15206 10092 15258
rect 9846 15204 9852 15206
rect 9908 15204 9932 15206
rect 9988 15204 10012 15206
rect 10068 15204 10092 15206
rect 10148 15204 10154 15206
rect 9846 15195 10154 15204
rect 7622 14716 7930 14725
rect 7622 14714 7628 14716
rect 7684 14714 7708 14716
rect 7764 14714 7788 14716
rect 7844 14714 7868 14716
rect 7924 14714 7930 14716
rect 7684 14662 7686 14714
rect 7866 14662 7868 14714
rect 7622 14660 7628 14662
rect 7684 14660 7708 14662
rect 7764 14660 7788 14662
rect 7844 14660 7868 14662
rect 7924 14660 7930 14662
rect 7622 14651 7930 14660
rect 5398 14172 5706 14181
rect 5398 14170 5404 14172
rect 5460 14170 5484 14172
rect 5540 14170 5564 14172
rect 5620 14170 5644 14172
rect 5700 14170 5706 14172
rect 5460 14118 5462 14170
rect 5642 14118 5644 14170
rect 5398 14116 5404 14118
rect 5460 14116 5484 14118
rect 5540 14116 5564 14118
rect 5620 14116 5644 14118
rect 5700 14116 5706 14118
rect 5398 14107 5706 14116
rect 9846 14172 10154 14181
rect 9846 14170 9852 14172
rect 9908 14170 9932 14172
rect 9988 14170 10012 14172
rect 10068 14170 10092 14172
rect 10148 14170 10154 14172
rect 9908 14118 9910 14170
rect 10090 14118 10092 14170
rect 9846 14116 9852 14118
rect 9908 14116 9932 14118
rect 9988 14116 10012 14118
rect 10068 14116 10092 14118
rect 10148 14116 10154 14118
rect 9846 14107 10154 14116
rect 7622 13628 7930 13637
rect 7622 13626 7628 13628
rect 7684 13626 7708 13628
rect 7764 13626 7788 13628
rect 7844 13626 7868 13628
rect 7924 13626 7930 13628
rect 7684 13574 7686 13626
rect 7866 13574 7868 13626
rect 7622 13572 7628 13574
rect 7684 13572 7708 13574
rect 7764 13572 7788 13574
rect 7844 13572 7868 13574
rect 7924 13572 7930 13574
rect 7622 13563 7930 13572
rect 5398 13084 5706 13093
rect 5398 13082 5404 13084
rect 5460 13082 5484 13084
rect 5540 13082 5564 13084
rect 5620 13082 5644 13084
rect 5700 13082 5706 13084
rect 5460 13030 5462 13082
rect 5642 13030 5644 13082
rect 5398 13028 5404 13030
rect 5460 13028 5484 13030
rect 5540 13028 5564 13030
rect 5620 13028 5644 13030
rect 5700 13028 5706 13030
rect 5398 13019 5706 13028
rect 9846 13084 10154 13093
rect 9846 13082 9852 13084
rect 9908 13082 9932 13084
rect 9988 13082 10012 13084
rect 10068 13082 10092 13084
rect 10148 13082 10154 13084
rect 9908 13030 9910 13082
rect 10090 13030 10092 13082
rect 9846 13028 9852 13030
rect 9908 13028 9932 13030
rect 9988 13028 10012 13030
rect 10068 13028 10092 13030
rect 10148 13028 10154 13030
rect 9846 13019 10154 13028
rect 7622 12540 7930 12549
rect 7622 12538 7628 12540
rect 7684 12538 7708 12540
rect 7764 12538 7788 12540
rect 7844 12538 7868 12540
rect 7924 12538 7930 12540
rect 7684 12486 7686 12538
rect 7866 12486 7868 12538
rect 7622 12484 7628 12486
rect 7684 12484 7708 12486
rect 7764 12484 7788 12486
rect 7844 12484 7868 12486
rect 7924 12484 7930 12486
rect 7622 12475 7930 12484
rect 10968 12096 11020 12102
rect 10968 12038 11020 12044
rect 5398 11996 5706 12005
rect 5398 11994 5404 11996
rect 5460 11994 5484 11996
rect 5540 11994 5564 11996
rect 5620 11994 5644 11996
rect 5700 11994 5706 11996
rect 5460 11942 5462 11994
rect 5642 11942 5644 11994
rect 5398 11940 5404 11942
rect 5460 11940 5484 11942
rect 5540 11940 5564 11942
rect 5620 11940 5644 11942
rect 5700 11940 5706 11942
rect 5398 11931 5706 11940
rect 9846 11996 10154 12005
rect 9846 11994 9852 11996
rect 9908 11994 9932 11996
rect 9988 11994 10012 11996
rect 10068 11994 10092 11996
rect 10148 11994 10154 11996
rect 9908 11942 9910 11994
rect 10090 11942 10092 11994
rect 9846 11940 9852 11942
rect 9908 11940 9932 11942
rect 9988 11940 10012 11942
rect 10068 11940 10092 11942
rect 10148 11940 10154 11942
rect 9846 11931 10154 11940
rect 10980 11898 11008 12038
rect 10968 11892 11020 11898
rect 10968 11834 11020 11840
rect 11532 11762 11560 16934
rect 12070 16892 12378 16901
rect 12070 16890 12076 16892
rect 12132 16890 12156 16892
rect 12212 16890 12236 16892
rect 12292 16890 12316 16892
rect 12372 16890 12378 16892
rect 12132 16838 12134 16890
rect 12314 16838 12316 16890
rect 12070 16836 12076 16838
rect 12132 16836 12156 16838
rect 12212 16836 12236 16838
rect 12292 16836 12316 16838
rect 12372 16836 12378 16838
rect 12070 16827 12378 16836
rect 16518 16892 16826 16901
rect 16518 16890 16524 16892
rect 16580 16890 16604 16892
rect 16660 16890 16684 16892
rect 16740 16890 16764 16892
rect 16820 16890 16826 16892
rect 16580 16838 16582 16890
rect 16762 16838 16764 16890
rect 16518 16836 16524 16838
rect 16580 16836 16604 16838
rect 16660 16836 16684 16838
rect 16740 16836 16764 16838
rect 16820 16836 16826 16838
rect 16518 16827 16826 16836
rect 14294 16348 14602 16357
rect 14294 16346 14300 16348
rect 14356 16346 14380 16348
rect 14436 16346 14460 16348
rect 14516 16346 14540 16348
rect 14596 16346 14602 16348
rect 14356 16294 14358 16346
rect 14538 16294 14540 16346
rect 14294 16292 14300 16294
rect 14356 16292 14380 16294
rect 14436 16292 14460 16294
rect 14516 16292 14540 16294
rect 14596 16292 14602 16294
rect 14294 16283 14602 16292
rect 12070 15804 12378 15813
rect 12070 15802 12076 15804
rect 12132 15802 12156 15804
rect 12212 15802 12236 15804
rect 12292 15802 12316 15804
rect 12372 15802 12378 15804
rect 12132 15750 12134 15802
rect 12314 15750 12316 15802
rect 12070 15748 12076 15750
rect 12132 15748 12156 15750
rect 12212 15748 12236 15750
rect 12292 15748 12316 15750
rect 12372 15748 12378 15750
rect 12070 15739 12378 15748
rect 16518 15804 16826 15813
rect 16518 15802 16524 15804
rect 16580 15802 16604 15804
rect 16660 15802 16684 15804
rect 16740 15802 16764 15804
rect 16820 15802 16826 15804
rect 16580 15750 16582 15802
rect 16762 15750 16764 15802
rect 16518 15748 16524 15750
rect 16580 15748 16604 15750
rect 16660 15748 16684 15750
rect 16740 15748 16764 15750
rect 16820 15748 16826 15750
rect 16518 15739 16826 15748
rect 14294 15260 14602 15269
rect 14294 15258 14300 15260
rect 14356 15258 14380 15260
rect 14436 15258 14460 15260
rect 14516 15258 14540 15260
rect 14596 15258 14602 15260
rect 14356 15206 14358 15258
rect 14538 15206 14540 15258
rect 14294 15204 14300 15206
rect 14356 15204 14380 15206
rect 14436 15204 14460 15206
rect 14516 15204 14540 15206
rect 14596 15204 14602 15206
rect 14294 15195 14602 15204
rect 12070 14716 12378 14725
rect 12070 14714 12076 14716
rect 12132 14714 12156 14716
rect 12212 14714 12236 14716
rect 12292 14714 12316 14716
rect 12372 14714 12378 14716
rect 12132 14662 12134 14714
rect 12314 14662 12316 14714
rect 12070 14660 12076 14662
rect 12132 14660 12156 14662
rect 12212 14660 12236 14662
rect 12292 14660 12316 14662
rect 12372 14660 12378 14662
rect 12070 14651 12378 14660
rect 16518 14716 16826 14725
rect 16518 14714 16524 14716
rect 16580 14714 16604 14716
rect 16660 14714 16684 14716
rect 16740 14714 16764 14716
rect 16820 14714 16826 14716
rect 16580 14662 16582 14714
rect 16762 14662 16764 14714
rect 16518 14660 16524 14662
rect 16580 14660 16604 14662
rect 16660 14660 16684 14662
rect 16740 14660 16764 14662
rect 16820 14660 16826 14662
rect 16518 14651 16826 14660
rect 14294 14172 14602 14181
rect 14294 14170 14300 14172
rect 14356 14170 14380 14172
rect 14436 14170 14460 14172
rect 14516 14170 14540 14172
rect 14596 14170 14602 14172
rect 14356 14118 14358 14170
rect 14538 14118 14540 14170
rect 14294 14116 14300 14118
rect 14356 14116 14380 14118
rect 14436 14116 14460 14118
rect 14516 14116 14540 14118
rect 14596 14116 14602 14118
rect 14294 14107 14602 14116
rect 12070 13628 12378 13637
rect 12070 13626 12076 13628
rect 12132 13626 12156 13628
rect 12212 13626 12236 13628
rect 12292 13626 12316 13628
rect 12372 13626 12378 13628
rect 12132 13574 12134 13626
rect 12314 13574 12316 13626
rect 12070 13572 12076 13574
rect 12132 13572 12156 13574
rect 12212 13572 12236 13574
rect 12292 13572 12316 13574
rect 12372 13572 12378 13574
rect 12070 13563 12378 13572
rect 16518 13628 16826 13637
rect 16518 13626 16524 13628
rect 16580 13626 16604 13628
rect 16660 13626 16684 13628
rect 16740 13626 16764 13628
rect 16820 13626 16826 13628
rect 16580 13574 16582 13626
rect 16762 13574 16764 13626
rect 16518 13572 16524 13574
rect 16580 13572 16604 13574
rect 16660 13572 16684 13574
rect 16740 13572 16764 13574
rect 16820 13572 16826 13574
rect 16518 13563 16826 13572
rect 14294 13084 14602 13093
rect 14294 13082 14300 13084
rect 14356 13082 14380 13084
rect 14436 13082 14460 13084
rect 14516 13082 14540 13084
rect 14596 13082 14602 13084
rect 14356 13030 14358 13082
rect 14538 13030 14540 13082
rect 14294 13028 14300 13030
rect 14356 13028 14380 13030
rect 14436 13028 14460 13030
rect 14516 13028 14540 13030
rect 14596 13028 14602 13030
rect 14294 13019 14602 13028
rect 12070 12540 12378 12549
rect 12070 12538 12076 12540
rect 12132 12538 12156 12540
rect 12212 12538 12236 12540
rect 12292 12538 12316 12540
rect 12372 12538 12378 12540
rect 12132 12486 12134 12538
rect 12314 12486 12316 12538
rect 12070 12484 12076 12486
rect 12132 12484 12156 12486
rect 12212 12484 12236 12486
rect 12292 12484 12316 12486
rect 12372 12484 12378 12486
rect 12070 12475 12378 12484
rect 16518 12540 16826 12549
rect 16518 12538 16524 12540
rect 16580 12538 16604 12540
rect 16660 12538 16684 12540
rect 16740 12538 16764 12540
rect 16820 12538 16826 12540
rect 16580 12486 16582 12538
rect 16762 12486 16764 12538
rect 16518 12484 16524 12486
rect 16580 12484 16604 12486
rect 16660 12484 16684 12486
rect 16740 12484 16764 12486
rect 16820 12484 16826 12486
rect 16518 12475 16826 12484
rect 12440 12300 12492 12306
rect 12440 12242 12492 12248
rect 11796 12096 11848 12102
rect 11796 12038 11848 12044
rect 11520 11756 11572 11762
rect 11520 11698 11572 11704
rect 4068 11552 4120 11558
rect 4068 11494 4120 11500
rect 3174 11452 3482 11461
rect 3174 11450 3180 11452
rect 3236 11450 3260 11452
rect 3316 11450 3340 11452
rect 3396 11450 3420 11452
rect 3476 11450 3482 11452
rect 3236 11398 3238 11450
rect 3418 11398 3420 11450
rect 3174 11396 3180 11398
rect 3236 11396 3260 11398
rect 3316 11396 3340 11398
rect 3396 11396 3420 11398
rect 3476 11396 3482 11398
rect 3174 11387 3482 11396
rect 7622 11452 7930 11461
rect 7622 11450 7628 11452
rect 7684 11450 7708 11452
rect 7764 11450 7788 11452
rect 7844 11450 7868 11452
rect 7924 11450 7930 11452
rect 7684 11398 7686 11450
rect 7866 11398 7868 11450
rect 7622 11396 7628 11398
rect 7684 11396 7708 11398
rect 7764 11396 7788 11398
rect 7844 11396 7868 11398
rect 7924 11396 7930 11398
rect 7622 11387 7930 11396
rect 10876 11280 10928 11286
rect 10876 11222 10928 11228
rect 20 11076 72 11082
rect 20 11018 72 11024
rect 32 800 60 11018
rect 5398 10908 5706 10917
rect 5398 10906 5404 10908
rect 5460 10906 5484 10908
rect 5540 10906 5564 10908
rect 5620 10906 5644 10908
rect 5700 10906 5706 10908
rect 5460 10854 5462 10906
rect 5642 10854 5644 10906
rect 5398 10852 5404 10854
rect 5460 10852 5484 10854
rect 5540 10852 5564 10854
rect 5620 10852 5644 10854
rect 5700 10852 5706 10854
rect 5398 10843 5706 10852
rect 9846 10908 10154 10917
rect 9846 10906 9852 10908
rect 9908 10906 9932 10908
rect 9988 10906 10012 10908
rect 10068 10906 10092 10908
rect 10148 10906 10154 10908
rect 9908 10854 9910 10906
rect 10090 10854 10092 10906
rect 9846 10852 9852 10854
rect 9908 10852 9932 10854
rect 9988 10852 10012 10854
rect 10068 10852 10092 10854
rect 10148 10852 10154 10854
rect 9846 10843 10154 10852
rect 10888 10674 10916 11222
rect 10416 10668 10468 10674
rect 10416 10610 10468 10616
rect 10876 10668 10928 10674
rect 10876 10610 10928 10616
rect 3174 10364 3482 10373
rect 3174 10362 3180 10364
rect 3236 10362 3260 10364
rect 3316 10362 3340 10364
rect 3396 10362 3420 10364
rect 3476 10362 3482 10364
rect 3236 10310 3238 10362
rect 3418 10310 3420 10362
rect 3174 10308 3180 10310
rect 3236 10308 3260 10310
rect 3316 10308 3340 10310
rect 3396 10308 3420 10310
rect 3476 10308 3482 10310
rect 3174 10299 3482 10308
rect 7622 10364 7930 10373
rect 7622 10362 7628 10364
rect 7684 10362 7708 10364
rect 7764 10362 7788 10364
rect 7844 10362 7868 10364
rect 7924 10362 7930 10364
rect 7684 10310 7686 10362
rect 7866 10310 7868 10362
rect 7622 10308 7628 10310
rect 7684 10308 7708 10310
rect 7764 10308 7788 10310
rect 7844 10308 7868 10310
rect 7924 10308 7930 10310
rect 7622 10299 7930 10308
rect 5398 9820 5706 9829
rect 5398 9818 5404 9820
rect 5460 9818 5484 9820
rect 5540 9818 5564 9820
rect 5620 9818 5644 9820
rect 5700 9818 5706 9820
rect 5460 9766 5462 9818
rect 5642 9766 5644 9818
rect 5398 9764 5404 9766
rect 5460 9764 5484 9766
rect 5540 9764 5564 9766
rect 5620 9764 5644 9766
rect 5700 9764 5706 9766
rect 5398 9755 5706 9764
rect 9846 9820 10154 9829
rect 9846 9818 9852 9820
rect 9908 9818 9932 9820
rect 9988 9818 10012 9820
rect 10068 9818 10092 9820
rect 10148 9818 10154 9820
rect 9908 9766 9910 9818
rect 10090 9766 10092 9818
rect 9846 9764 9852 9766
rect 9908 9764 9932 9766
rect 9988 9764 10012 9766
rect 10068 9764 10092 9766
rect 10148 9764 10154 9766
rect 9846 9755 10154 9764
rect 3174 9276 3482 9285
rect 3174 9274 3180 9276
rect 3236 9274 3260 9276
rect 3316 9274 3340 9276
rect 3396 9274 3420 9276
rect 3476 9274 3482 9276
rect 3236 9222 3238 9274
rect 3418 9222 3420 9274
rect 3174 9220 3180 9222
rect 3236 9220 3260 9222
rect 3316 9220 3340 9222
rect 3396 9220 3420 9222
rect 3476 9220 3482 9222
rect 3174 9211 3482 9220
rect 7622 9276 7930 9285
rect 7622 9274 7628 9276
rect 7684 9274 7708 9276
rect 7764 9274 7788 9276
rect 7844 9274 7868 9276
rect 7924 9274 7930 9276
rect 7684 9222 7686 9274
rect 7866 9222 7868 9274
rect 7622 9220 7628 9222
rect 7684 9220 7708 9222
rect 7764 9220 7788 9222
rect 7844 9220 7868 9222
rect 7924 9220 7930 9222
rect 7622 9211 7930 9220
rect 5398 8732 5706 8741
rect 5398 8730 5404 8732
rect 5460 8730 5484 8732
rect 5540 8730 5564 8732
rect 5620 8730 5644 8732
rect 5700 8730 5706 8732
rect 5460 8678 5462 8730
rect 5642 8678 5644 8730
rect 5398 8676 5404 8678
rect 5460 8676 5484 8678
rect 5540 8676 5564 8678
rect 5620 8676 5644 8678
rect 5700 8676 5706 8678
rect 5398 8667 5706 8676
rect 9846 8732 10154 8741
rect 9846 8730 9852 8732
rect 9908 8730 9932 8732
rect 9988 8730 10012 8732
rect 10068 8730 10092 8732
rect 10148 8730 10154 8732
rect 9908 8678 9910 8730
rect 10090 8678 10092 8730
rect 9846 8676 9852 8678
rect 9908 8676 9932 8678
rect 9988 8676 10012 8678
rect 10068 8676 10092 8678
rect 10148 8676 10154 8678
rect 9846 8667 10154 8676
rect 3174 8188 3482 8197
rect 3174 8186 3180 8188
rect 3236 8186 3260 8188
rect 3316 8186 3340 8188
rect 3396 8186 3420 8188
rect 3476 8186 3482 8188
rect 3236 8134 3238 8186
rect 3418 8134 3420 8186
rect 3174 8132 3180 8134
rect 3236 8132 3260 8134
rect 3316 8132 3340 8134
rect 3396 8132 3420 8134
rect 3476 8132 3482 8134
rect 3174 8123 3482 8132
rect 7622 8188 7930 8197
rect 7622 8186 7628 8188
rect 7684 8186 7708 8188
rect 7764 8186 7788 8188
rect 7844 8186 7868 8188
rect 7924 8186 7930 8188
rect 7684 8134 7686 8186
rect 7866 8134 7868 8186
rect 7622 8132 7628 8134
rect 7684 8132 7708 8134
rect 7764 8132 7788 8134
rect 7844 8132 7868 8134
rect 7924 8132 7930 8134
rect 7622 8123 7930 8132
rect 10428 7886 10456 10610
rect 11808 10062 11836 12038
rect 12452 11898 12480 12242
rect 12808 12232 12860 12238
rect 12808 12174 12860 12180
rect 12440 11892 12492 11898
rect 12440 11834 12492 11840
rect 12820 11558 12848 12174
rect 14294 11996 14602 12005
rect 14294 11994 14300 11996
rect 14356 11994 14380 11996
rect 14436 11994 14460 11996
rect 14516 11994 14540 11996
rect 14596 11994 14602 11996
rect 14356 11942 14358 11994
rect 14538 11942 14540 11994
rect 14294 11940 14300 11942
rect 14356 11940 14380 11942
rect 14436 11940 14460 11942
rect 14516 11940 14540 11942
rect 14596 11940 14602 11942
rect 14294 11931 14602 11940
rect 12900 11892 12952 11898
rect 12900 11834 12952 11840
rect 12716 11552 12768 11558
rect 12716 11494 12768 11500
rect 12808 11552 12860 11558
rect 12808 11494 12860 11500
rect 12070 11452 12378 11461
rect 12070 11450 12076 11452
rect 12132 11450 12156 11452
rect 12212 11450 12236 11452
rect 12292 11450 12316 11452
rect 12372 11450 12378 11452
rect 12132 11398 12134 11450
rect 12314 11398 12316 11450
rect 12070 11396 12076 11398
rect 12132 11396 12156 11398
rect 12212 11396 12236 11398
rect 12292 11396 12316 11398
rect 12372 11396 12378 11398
rect 12070 11387 12378 11396
rect 12728 11150 12756 11494
rect 12716 11144 12768 11150
rect 12716 11086 12768 11092
rect 12440 11076 12492 11082
rect 12440 11018 12492 11024
rect 12452 10742 12480 11018
rect 12440 10736 12492 10742
rect 12440 10678 12492 10684
rect 12070 10364 12378 10373
rect 12070 10362 12076 10364
rect 12132 10362 12156 10364
rect 12212 10362 12236 10364
rect 12292 10362 12316 10364
rect 12372 10362 12378 10364
rect 12132 10310 12134 10362
rect 12314 10310 12316 10362
rect 12070 10308 12076 10310
rect 12132 10308 12156 10310
rect 12212 10308 12236 10310
rect 12292 10308 12316 10310
rect 12372 10308 12378 10310
rect 12070 10299 12378 10308
rect 12912 10266 12940 11834
rect 18144 11756 18196 11762
rect 18144 11698 18196 11704
rect 18156 11665 18184 11698
rect 18142 11656 18198 11665
rect 18142 11591 18198 11600
rect 14556 11552 14608 11558
rect 14556 11494 14608 11500
rect 14568 11150 14596 11494
rect 16518 11452 16826 11461
rect 16518 11450 16524 11452
rect 16580 11450 16604 11452
rect 16660 11450 16684 11452
rect 16740 11450 16764 11452
rect 16820 11450 16826 11452
rect 16580 11398 16582 11450
rect 16762 11398 16764 11450
rect 16518 11396 16524 11398
rect 16580 11396 16604 11398
rect 16660 11396 16684 11398
rect 16740 11396 16764 11398
rect 16820 11396 16826 11398
rect 16518 11387 16826 11396
rect 14556 11144 14608 11150
rect 14556 11086 14608 11092
rect 13820 11008 13872 11014
rect 13820 10950 13872 10956
rect 15568 11008 15620 11014
rect 15568 10950 15620 10956
rect 13832 10810 13860 10950
rect 14294 10908 14602 10917
rect 14294 10906 14300 10908
rect 14356 10906 14380 10908
rect 14436 10906 14460 10908
rect 14516 10906 14540 10908
rect 14596 10906 14602 10908
rect 14356 10854 14358 10906
rect 14538 10854 14540 10906
rect 14294 10852 14300 10854
rect 14356 10852 14380 10854
rect 14436 10852 14460 10854
rect 14516 10852 14540 10854
rect 14596 10852 14602 10854
rect 14294 10843 14602 10852
rect 13820 10804 13872 10810
rect 13820 10746 13872 10752
rect 12900 10260 12952 10266
rect 12900 10202 12952 10208
rect 11612 10056 11664 10062
rect 11612 9998 11664 10004
rect 11796 10056 11848 10062
rect 11796 9998 11848 10004
rect 11624 9674 11652 9998
rect 14294 9820 14602 9829
rect 14294 9818 14300 9820
rect 14356 9818 14380 9820
rect 14436 9818 14460 9820
rect 14516 9818 14540 9820
rect 14596 9818 14602 9820
rect 14356 9766 14358 9818
rect 14538 9766 14540 9818
rect 14294 9764 14300 9766
rect 14356 9764 14380 9766
rect 14436 9764 14460 9766
rect 14516 9764 14540 9766
rect 14596 9764 14602 9766
rect 14294 9755 14602 9764
rect 11624 9646 11744 9674
rect 11716 8090 11744 9646
rect 12070 9276 12378 9285
rect 12070 9274 12076 9276
rect 12132 9274 12156 9276
rect 12212 9274 12236 9276
rect 12292 9274 12316 9276
rect 12372 9274 12378 9276
rect 12132 9222 12134 9274
rect 12314 9222 12316 9274
rect 12070 9220 12076 9222
rect 12132 9220 12156 9222
rect 12212 9220 12236 9222
rect 12292 9220 12316 9222
rect 12372 9220 12378 9222
rect 12070 9211 12378 9220
rect 14294 8732 14602 8741
rect 14294 8730 14300 8732
rect 14356 8730 14380 8732
rect 14436 8730 14460 8732
rect 14516 8730 14540 8732
rect 14596 8730 14602 8732
rect 14356 8678 14358 8730
rect 14538 8678 14540 8730
rect 14294 8676 14300 8678
rect 14356 8676 14380 8678
rect 14436 8676 14460 8678
rect 14516 8676 14540 8678
rect 14596 8676 14602 8678
rect 14294 8667 14602 8676
rect 12070 8188 12378 8197
rect 12070 8186 12076 8188
rect 12132 8186 12156 8188
rect 12212 8186 12236 8188
rect 12292 8186 12316 8188
rect 12372 8186 12378 8188
rect 12132 8134 12134 8186
rect 12314 8134 12316 8186
rect 12070 8132 12076 8134
rect 12132 8132 12156 8134
rect 12212 8132 12236 8134
rect 12292 8132 12316 8134
rect 12372 8132 12378 8134
rect 12070 8123 12378 8132
rect 11704 8084 11756 8090
rect 11704 8026 11756 8032
rect 10416 7880 10468 7886
rect 10416 7822 10468 7828
rect 5398 7644 5706 7653
rect 5398 7642 5404 7644
rect 5460 7642 5484 7644
rect 5540 7642 5564 7644
rect 5620 7642 5644 7644
rect 5700 7642 5706 7644
rect 5460 7590 5462 7642
rect 5642 7590 5644 7642
rect 5398 7588 5404 7590
rect 5460 7588 5484 7590
rect 5540 7588 5564 7590
rect 5620 7588 5644 7590
rect 5700 7588 5706 7590
rect 5398 7579 5706 7588
rect 9846 7644 10154 7653
rect 9846 7642 9852 7644
rect 9908 7642 9932 7644
rect 9988 7642 10012 7644
rect 10068 7642 10092 7644
rect 10148 7642 10154 7644
rect 9908 7590 9910 7642
rect 10090 7590 10092 7642
rect 9846 7588 9852 7590
rect 9908 7588 9932 7590
rect 9988 7588 10012 7590
rect 10068 7588 10092 7590
rect 10148 7588 10154 7590
rect 9846 7579 10154 7588
rect 14294 7644 14602 7653
rect 14294 7642 14300 7644
rect 14356 7642 14380 7644
rect 14436 7642 14460 7644
rect 14516 7642 14540 7644
rect 14596 7642 14602 7644
rect 14356 7590 14358 7642
rect 14538 7590 14540 7642
rect 14294 7588 14300 7590
rect 14356 7588 14380 7590
rect 14436 7588 14460 7590
rect 14516 7588 14540 7590
rect 14596 7588 14602 7590
rect 14294 7579 14602 7588
rect 3174 7100 3482 7109
rect 3174 7098 3180 7100
rect 3236 7098 3260 7100
rect 3316 7098 3340 7100
rect 3396 7098 3420 7100
rect 3476 7098 3482 7100
rect 3236 7046 3238 7098
rect 3418 7046 3420 7098
rect 3174 7044 3180 7046
rect 3236 7044 3260 7046
rect 3316 7044 3340 7046
rect 3396 7044 3420 7046
rect 3476 7044 3482 7046
rect 3174 7035 3482 7044
rect 7622 7100 7930 7109
rect 7622 7098 7628 7100
rect 7684 7098 7708 7100
rect 7764 7098 7788 7100
rect 7844 7098 7868 7100
rect 7924 7098 7930 7100
rect 7684 7046 7686 7098
rect 7866 7046 7868 7098
rect 7622 7044 7628 7046
rect 7684 7044 7708 7046
rect 7764 7044 7788 7046
rect 7844 7044 7868 7046
rect 7924 7044 7930 7046
rect 7622 7035 7930 7044
rect 12070 7100 12378 7109
rect 12070 7098 12076 7100
rect 12132 7098 12156 7100
rect 12212 7098 12236 7100
rect 12292 7098 12316 7100
rect 12372 7098 12378 7100
rect 12132 7046 12134 7098
rect 12314 7046 12316 7098
rect 12070 7044 12076 7046
rect 12132 7044 12156 7046
rect 12212 7044 12236 7046
rect 12292 7044 12316 7046
rect 12372 7044 12378 7046
rect 12070 7035 12378 7044
rect 5398 6556 5706 6565
rect 5398 6554 5404 6556
rect 5460 6554 5484 6556
rect 5540 6554 5564 6556
rect 5620 6554 5644 6556
rect 5700 6554 5706 6556
rect 5460 6502 5462 6554
rect 5642 6502 5644 6554
rect 5398 6500 5404 6502
rect 5460 6500 5484 6502
rect 5540 6500 5564 6502
rect 5620 6500 5644 6502
rect 5700 6500 5706 6502
rect 5398 6491 5706 6500
rect 9846 6556 10154 6565
rect 9846 6554 9852 6556
rect 9908 6554 9932 6556
rect 9988 6554 10012 6556
rect 10068 6554 10092 6556
rect 10148 6554 10154 6556
rect 9908 6502 9910 6554
rect 10090 6502 10092 6554
rect 9846 6500 9852 6502
rect 9908 6500 9932 6502
rect 9988 6500 10012 6502
rect 10068 6500 10092 6502
rect 10148 6500 10154 6502
rect 9846 6491 10154 6500
rect 14294 6556 14602 6565
rect 14294 6554 14300 6556
rect 14356 6554 14380 6556
rect 14436 6554 14460 6556
rect 14516 6554 14540 6556
rect 14596 6554 14602 6556
rect 14356 6502 14358 6554
rect 14538 6502 14540 6554
rect 14294 6500 14300 6502
rect 14356 6500 14380 6502
rect 14436 6500 14460 6502
rect 14516 6500 14540 6502
rect 14596 6500 14602 6502
rect 14294 6491 14602 6500
rect 3174 6012 3482 6021
rect 3174 6010 3180 6012
rect 3236 6010 3260 6012
rect 3316 6010 3340 6012
rect 3396 6010 3420 6012
rect 3476 6010 3482 6012
rect 3236 5958 3238 6010
rect 3418 5958 3420 6010
rect 3174 5956 3180 5958
rect 3236 5956 3260 5958
rect 3316 5956 3340 5958
rect 3396 5956 3420 5958
rect 3476 5956 3482 5958
rect 3174 5947 3482 5956
rect 7622 6012 7930 6021
rect 7622 6010 7628 6012
rect 7684 6010 7708 6012
rect 7764 6010 7788 6012
rect 7844 6010 7868 6012
rect 7924 6010 7930 6012
rect 7684 5958 7686 6010
rect 7866 5958 7868 6010
rect 7622 5956 7628 5958
rect 7684 5956 7708 5958
rect 7764 5956 7788 5958
rect 7844 5956 7868 5958
rect 7924 5956 7930 5958
rect 7622 5947 7930 5956
rect 12070 6012 12378 6021
rect 12070 6010 12076 6012
rect 12132 6010 12156 6012
rect 12212 6010 12236 6012
rect 12292 6010 12316 6012
rect 12372 6010 12378 6012
rect 12132 5958 12134 6010
rect 12314 5958 12316 6010
rect 12070 5956 12076 5958
rect 12132 5956 12156 5958
rect 12212 5956 12236 5958
rect 12292 5956 12316 5958
rect 12372 5956 12378 5958
rect 12070 5947 12378 5956
rect 5398 5468 5706 5477
rect 5398 5466 5404 5468
rect 5460 5466 5484 5468
rect 5540 5466 5564 5468
rect 5620 5466 5644 5468
rect 5700 5466 5706 5468
rect 5460 5414 5462 5466
rect 5642 5414 5644 5466
rect 5398 5412 5404 5414
rect 5460 5412 5484 5414
rect 5540 5412 5564 5414
rect 5620 5412 5644 5414
rect 5700 5412 5706 5414
rect 5398 5403 5706 5412
rect 9846 5468 10154 5477
rect 9846 5466 9852 5468
rect 9908 5466 9932 5468
rect 9988 5466 10012 5468
rect 10068 5466 10092 5468
rect 10148 5466 10154 5468
rect 9908 5414 9910 5466
rect 10090 5414 10092 5466
rect 9846 5412 9852 5414
rect 9908 5412 9932 5414
rect 9988 5412 10012 5414
rect 10068 5412 10092 5414
rect 10148 5412 10154 5414
rect 9846 5403 10154 5412
rect 14294 5468 14602 5477
rect 14294 5466 14300 5468
rect 14356 5466 14380 5468
rect 14436 5466 14460 5468
rect 14516 5466 14540 5468
rect 14596 5466 14602 5468
rect 14356 5414 14358 5466
rect 14538 5414 14540 5466
rect 14294 5412 14300 5414
rect 14356 5412 14380 5414
rect 14436 5412 14460 5414
rect 14516 5412 14540 5414
rect 14596 5412 14602 5414
rect 14294 5403 14602 5412
rect 3174 4924 3482 4933
rect 3174 4922 3180 4924
rect 3236 4922 3260 4924
rect 3316 4922 3340 4924
rect 3396 4922 3420 4924
rect 3476 4922 3482 4924
rect 3236 4870 3238 4922
rect 3418 4870 3420 4922
rect 3174 4868 3180 4870
rect 3236 4868 3260 4870
rect 3316 4868 3340 4870
rect 3396 4868 3420 4870
rect 3476 4868 3482 4870
rect 3174 4859 3482 4868
rect 7622 4924 7930 4933
rect 7622 4922 7628 4924
rect 7684 4922 7708 4924
rect 7764 4922 7788 4924
rect 7844 4922 7868 4924
rect 7924 4922 7930 4924
rect 7684 4870 7686 4922
rect 7866 4870 7868 4922
rect 7622 4868 7628 4870
rect 7684 4868 7708 4870
rect 7764 4868 7788 4870
rect 7844 4868 7868 4870
rect 7924 4868 7930 4870
rect 7622 4859 7930 4868
rect 12070 4924 12378 4933
rect 12070 4922 12076 4924
rect 12132 4922 12156 4924
rect 12212 4922 12236 4924
rect 12292 4922 12316 4924
rect 12372 4922 12378 4924
rect 12132 4870 12134 4922
rect 12314 4870 12316 4922
rect 12070 4868 12076 4870
rect 12132 4868 12156 4870
rect 12212 4868 12236 4870
rect 12292 4868 12316 4870
rect 12372 4868 12378 4870
rect 12070 4859 12378 4868
rect 5398 4380 5706 4389
rect 5398 4378 5404 4380
rect 5460 4378 5484 4380
rect 5540 4378 5564 4380
rect 5620 4378 5644 4380
rect 5700 4378 5706 4380
rect 5460 4326 5462 4378
rect 5642 4326 5644 4378
rect 5398 4324 5404 4326
rect 5460 4324 5484 4326
rect 5540 4324 5564 4326
rect 5620 4324 5644 4326
rect 5700 4324 5706 4326
rect 5398 4315 5706 4324
rect 9846 4380 10154 4389
rect 9846 4378 9852 4380
rect 9908 4378 9932 4380
rect 9988 4378 10012 4380
rect 10068 4378 10092 4380
rect 10148 4378 10154 4380
rect 9908 4326 9910 4378
rect 10090 4326 10092 4378
rect 9846 4324 9852 4326
rect 9908 4324 9932 4326
rect 9988 4324 10012 4326
rect 10068 4324 10092 4326
rect 10148 4324 10154 4326
rect 9846 4315 10154 4324
rect 14294 4380 14602 4389
rect 14294 4378 14300 4380
rect 14356 4378 14380 4380
rect 14436 4378 14460 4380
rect 14516 4378 14540 4380
rect 14596 4378 14602 4380
rect 14356 4326 14358 4378
rect 14538 4326 14540 4378
rect 14294 4324 14300 4326
rect 14356 4324 14380 4326
rect 14436 4324 14460 4326
rect 14516 4324 14540 4326
rect 14596 4324 14602 4326
rect 14294 4315 14602 4324
rect 3174 3836 3482 3845
rect 3174 3834 3180 3836
rect 3236 3834 3260 3836
rect 3316 3834 3340 3836
rect 3396 3834 3420 3836
rect 3476 3834 3482 3836
rect 3236 3782 3238 3834
rect 3418 3782 3420 3834
rect 3174 3780 3180 3782
rect 3236 3780 3260 3782
rect 3316 3780 3340 3782
rect 3396 3780 3420 3782
rect 3476 3780 3482 3782
rect 3174 3771 3482 3780
rect 7622 3836 7930 3845
rect 7622 3834 7628 3836
rect 7684 3834 7708 3836
rect 7764 3834 7788 3836
rect 7844 3834 7868 3836
rect 7924 3834 7930 3836
rect 7684 3782 7686 3834
rect 7866 3782 7868 3834
rect 7622 3780 7628 3782
rect 7684 3780 7708 3782
rect 7764 3780 7788 3782
rect 7844 3780 7868 3782
rect 7924 3780 7930 3782
rect 7622 3771 7930 3780
rect 12070 3836 12378 3845
rect 12070 3834 12076 3836
rect 12132 3834 12156 3836
rect 12212 3834 12236 3836
rect 12292 3834 12316 3836
rect 12372 3834 12378 3836
rect 12132 3782 12134 3834
rect 12314 3782 12316 3834
rect 12070 3780 12076 3782
rect 12132 3780 12156 3782
rect 12212 3780 12236 3782
rect 12292 3780 12316 3782
rect 12372 3780 12378 3782
rect 12070 3771 12378 3780
rect 5398 3292 5706 3301
rect 5398 3290 5404 3292
rect 5460 3290 5484 3292
rect 5540 3290 5564 3292
rect 5620 3290 5644 3292
rect 5700 3290 5706 3292
rect 5460 3238 5462 3290
rect 5642 3238 5644 3290
rect 5398 3236 5404 3238
rect 5460 3236 5484 3238
rect 5540 3236 5564 3238
rect 5620 3236 5644 3238
rect 5700 3236 5706 3238
rect 5398 3227 5706 3236
rect 9846 3292 10154 3301
rect 9846 3290 9852 3292
rect 9908 3290 9932 3292
rect 9988 3290 10012 3292
rect 10068 3290 10092 3292
rect 10148 3290 10154 3292
rect 9908 3238 9910 3290
rect 10090 3238 10092 3290
rect 9846 3236 9852 3238
rect 9908 3236 9932 3238
rect 9988 3236 10012 3238
rect 10068 3236 10092 3238
rect 10148 3236 10154 3238
rect 9846 3227 10154 3236
rect 14294 3292 14602 3301
rect 14294 3290 14300 3292
rect 14356 3290 14380 3292
rect 14436 3290 14460 3292
rect 14516 3290 14540 3292
rect 14596 3290 14602 3292
rect 14356 3238 14358 3290
rect 14538 3238 14540 3290
rect 14294 3236 14300 3238
rect 14356 3236 14380 3238
rect 14436 3236 14460 3238
rect 14516 3236 14540 3238
rect 14596 3236 14602 3238
rect 14294 3227 14602 3236
rect 3174 2748 3482 2757
rect 3174 2746 3180 2748
rect 3236 2746 3260 2748
rect 3316 2746 3340 2748
rect 3396 2746 3420 2748
rect 3476 2746 3482 2748
rect 3236 2694 3238 2746
rect 3418 2694 3420 2746
rect 3174 2692 3180 2694
rect 3236 2692 3260 2694
rect 3316 2692 3340 2694
rect 3396 2692 3420 2694
rect 3476 2692 3482 2694
rect 3174 2683 3482 2692
rect 7622 2748 7930 2757
rect 7622 2746 7628 2748
rect 7684 2746 7708 2748
rect 7764 2746 7788 2748
rect 7844 2746 7868 2748
rect 7924 2746 7930 2748
rect 7684 2694 7686 2746
rect 7866 2694 7868 2746
rect 7622 2692 7628 2694
rect 7684 2692 7708 2694
rect 7764 2692 7788 2694
rect 7844 2692 7868 2694
rect 7924 2692 7930 2694
rect 7622 2683 7930 2692
rect 12070 2748 12378 2757
rect 12070 2746 12076 2748
rect 12132 2746 12156 2748
rect 12212 2746 12236 2748
rect 12292 2746 12316 2748
rect 12372 2746 12378 2748
rect 12132 2694 12134 2746
rect 12314 2694 12316 2746
rect 12070 2692 12076 2694
rect 12132 2692 12156 2694
rect 12212 2692 12236 2694
rect 12292 2692 12316 2694
rect 12372 2692 12378 2694
rect 12070 2683 12378 2692
rect 15580 2446 15608 10950
rect 16518 10364 16826 10373
rect 16518 10362 16524 10364
rect 16580 10362 16604 10364
rect 16660 10362 16684 10364
rect 16740 10362 16764 10364
rect 16820 10362 16826 10364
rect 16580 10310 16582 10362
rect 16762 10310 16764 10362
rect 16518 10308 16524 10310
rect 16580 10308 16604 10310
rect 16660 10308 16684 10310
rect 16740 10308 16764 10310
rect 16820 10308 16826 10310
rect 16518 10299 16826 10308
rect 16518 9276 16826 9285
rect 16518 9274 16524 9276
rect 16580 9274 16604 9276
rect 16660 9274 16684 9276
rect 16740 9274 16764 9276
rect 16820 9274 16826 9276
rect 16580 9222 16582 9274
rect 16762 9222 16764 9274
rect 16518 9220 16524 9222
rect 16580 9220 16604 9222
rect 16660 9220 16684 9222
rect 16740 9220 16764 9222
rect 16820 9220 16826 9222
rect 16518 9211 16826 9220
rect 16518 8188 16826 8197
rect 16518 8186 16524 8188
rect 16580 8186 16604 8188
rect 16660 8186 16684 8188
rect 16740 8186 16764 8188
rect 16820 8186 16826 8188
rect 16580 8134 16582 8186
rect 16762 8134 16764 8186
rect 16518 8132 16524 8134
rect 16580 8132 16604 8134
rect 16660 8132 16684 8134
rect 16740 8132 16764 8134
rect 16820 8132 16826 8134
rect 16518 8123 16826 8132
rect 16518 7100 16826 7109
rect 16518 7098 16524 7100
rect 16580 7098 16604 7100
rect 16660 7098 16684 7100
rect 16740 7098 16764 7100
rect 16820 7098 16826 7100
rect 16580 7046 16582 7098
rect 16762 7046 16764 7098
rect 16518 7044 16524 7046
rect 16580 7044 16604 7046
rect 16660 7044 16684 7046
rect 16740 7044 16764 7046
rect 16820 7044 16826 7046
rect 16518 7035 16826 7044
rect 16518 6012 16826 6021
rect 16518 6010 16524 6012
rect 16580 6010 16604 6012
rect 16660 6010 16684 6012
rect 16740 6010 16764 6012
rect 16820 6010 16826 6012
rect 16580 5958 16582 6010
rect 16762 5958 16764 6010
rect 16518 5956 16524 5958
rect 16580 5956 16604 5958
rect 16660 5956 16684 5958
rect 16740 5956 16764 5958
rect 16820 5956 16826 5958
rect 16518 5947 16826 5956
rect 16518 4924 16826 4933
rect 16518 4922 16524 4924
rect 16580 4922 16604 4924
rect 16660 4922 16684 4924
rect 16740 4922 16764 4924
rect 16820 4922 16826 4924
rect 16580 4870 16582 4922
rect 16762 4870 16764 4922
rect 16518 4868 16524 4870
rect 16580 4868 16604 4870
rect 16660 4868 16684 4870
rect 16740 4868 16764 4870
rect 16820 4868 16826 4870
rect 16518 4859 16826 4868
rect 16518 3836 16826 3845
rect 16518 3834 16524 3836
rect 16580 3834 16604 3836
rect 16660 3834 16684 3836
rect 16740 3834 16764 3836
rect 16820 3834 16826 3836
rect 16580 3782 16582 3834
rect 16762 3782 16764 3834
rect 16518 3780 16524 3782
rect 16580 3780 16604 3782
rect 16660 3780 16684 3782
rect 16740 3780 16764 3782
rect 16820 3780 16826 3782
rect 16518 3771 16826 3780
rect 16518 2748 16826 2757
rect 16518 2746 16524 2748
rect 16580 2746 16604 2748
rect 16660 2746 16684 2748
rect 16740 2746 16764 2748
rect 16820 2746 16826 2748
rect 16580 2694 16582 2746
rect 16762 2694 16764 2746
rect 16518 2692 16524 2694
rect 16580 2692 16604 2694
rect 16660 2692 16684 2694
rect 16740 2692 16764 2694
rect 16820 2692 16826 2694
rect 16518 2683 16826 2692
rect 15568 2440 15620 2446
rect 15568 2382 15620 2388
rect 15476 2304 15528 2310
rect 15476 2246 15528 2252
rect 5398 2204 5706 2213
rect 5398 2202 5404 2204
rect 5460 2202 5484 2204
rect 5540 2202 5564 2204
rect 5620 2202 5644 2204
rect 5700 2202 5706 2204
rect 5460 2150 5462 2202
rect 5642 2150 5644 2202
rect 5398 2148 5404 2150
rect 5460 2148 5484 2150
rect 5540 2148 5564 2150
rect 5620 2148 5644 2150
rect 5700 2148 5706 2150
rect 5398 2139 5706 2148
rect 9846 2204 10154 2213
rect 9846 2202 9852 2204
rect 9908 2202 9932 2204
rect 9988 2202 10012 2204
rect 10068 2202 10092 2204
rect 10148 2202 10154 2204
rect 9908 2150 9910 2202
rect 10090 2150 10092 2202
rect 9846 2148 9852 2150
rect 9908 2148 9932 2150
rect 9988 2148 10012 2150
rect 10068 2148 10092 2150
rect 10148 2148 10154 2150
rect 9846 2139 10154 2148
rect 14294 2204 14602 2213
rect 14294 2202 14300 2204
rect 14356 2202 14380 2204
rect 14436 2202 14460 2204
rect 14516 2202 14540 2204
rect 14596 2202 14602 2204
rect 14356 2150 14358 2202
rect 14538 2150 14540 2202
rect 14294 2148 14300 2150
rect 14356 2148 14380 2150
rect 14436 2148 14460 2150
rect 14516 2148 14540 2150
rect 14596 2148 14602 2150
rect 14294 2139 14602 2148
rect 15488 800 15516 2246
rect 18 0 74 800
rect 15474 0 15530 800
<< via2 >>
rect 5404 17434 5460 17436
rect 5484 17434 5540 17436
rect 5564 17434 5620 17436
rect 5644 17434 5700 17436
rect 5404 17382 5450 17434
rect 5450 17382 5460 17434
rect 5484 17382 5514 17434
rect 5514 17382 5526 17434
rect 5526 17382 5540 17434
rect 5564 17382 5578 17434
rect 5578 17382 5590 17434
rect 5590 17382 5620 17434
rect 5644 17382 5654 17434
rect 5654 17382 5700 17434
rect 5404 17380 5460 17382
rect 5484 17380 5540 17382
rect 5564 17380 5620 17382
rect 5644 17380 5700 17382
rect 9852 17434 9908 17436
rect 9932 17434 9988 17436
rect 10012 17434 10068 17436
rect 10092 17434 10148 17436
rect 9852 17382 9898 17434
rect 9898 17382 9908 17434
rect 9932 17382 9962 17434
rect 9962 17382 9974 17434
rect 9974 17382 9988 17434
rect 10012 17382 10026 17434
rect 10026 17382 10038 17434
rect 10038 17382 10068 17434
rect 10092 17382 10102 17434
rect 10102 17382 10148 17434
rect 9852 17380 9908 17382
rect 9932 17380 9988 17382
rect 10012 17380 10068 17382
rect 10092 17380 10148 17382
rect 14300 17434 14356 17436
rect 14380 17434 14436 17436
rect 14460 17434 14516 17436
rect 14540 17434 14596 17436
rect 14300 17382 14346 17434
rect 14346 17382 14356 17434
rect 14380 17382 14410 17434
rect 14410 17382 14422 17434
rect 14422 17382 14436 17434
rect 14460 17382 14474 17434
rect 14474 17382 14486 17434
rect 14486 17382 14516 17434
rect 14540 17382 14550 17434
rect 14550 17382 14596 17434
rect 14300 17380 14356 17382
rect 14380 17380 14436 17382
rect 14460 17380 14516 17382
rect 14540 17380 14596 17382
rect 3180 16890 3236 16892
rect 3260 16890 3316 16892
rect 3340 16890 3396 16892
rect 3420 16890 3476 16892
rect 3180 16838 3226 16890
rect 3226 16838 3236 16890
rect 3260 16838 3290 16890
rect 3290 16838 3302 16890
rect 3302 16838 3316 16890
rect 3340 16838 3354 16890
rect 3354 16838 3366 16890
rect 3366 16838 3396 16890
rect 3420 16838 3430 16890
rect 3430 16838 3476 16890
rect 3180 16836 3236 16838
rect 3260 16836 3316 16838
rect 3340 16836 3396 16838
rect 3420 16836 3476 16838
rect 7628 16890 7684 16892
rect 7708 16890 7764 16892
rect 7788 16890 7844 16892
rect 7868 16890 7924 16892
rect 7628 16838 7674 16890
rect 7674 16838 7684 16890
rect 7708 16838 7738 16890
rect 7738 16838 7750 16890
rect 7750 16838 7764 16890
rect 7788 16838 7802 16890
rect 7802 16838 7814 16890
rect 7814 16838 7844 16890
rect 7868 16838 7878 16890
rect 7878 16838 7924 16890
rect 7628 16836 7684 16838
rect 7708 16836 7764 16838
rect 7788 16836 7844 16838
rect 7868 16836 7924 16838
rect 1398 16360 1454 16416
rect 3180 15802 3236 15804
rect 3260 15802 3316 15804
rect 3340 15802 3396 15804
rect 3420 15802 3476 15804
rect 3180 15750 3226 15802
rect 3226 15750 3236 15802
rect 3260 15750 3290 15802
rect 3290 15750 3302 15802
rect 3302 15750 3316 15802
rect 3340 15750 3354 15802
rect 3354 15750 3366 15802
rect 3366 15750 3396 15802
rect 3420 15750 3430 15802
rect 3430 15750 3476 15802
rect 3180 15748 3236 15750
rect 3260 15748 3316 15750
rect 3340 15748 3396 15750
rect 3420 15748 3476 15750
rect 3180 14714 3236 14716
rect 3260 14714 3316 14716
rect 3340 14714 3396 14716
rect 3420 14714 3476 14716
rect 3180 14662 3226 14714
rect 3226 14662 3236 14714
rect 3260 14662 3290 14714
rect 3290 14662 3302 14714
rect 3302 14662 3316 14714
rect 3340 14662 3354 14714
rect 3354 14662 3366 14714
rect 3366 14662 3396 14714
rect 3420 14662 3430 14714
rect 3430 14662 3476 14714
rect 3180 14660 3236 14662
rect 3260 14660 3316 14662
rect 3340 14660 3396 14662
rect 3420 14660 3476 14662
rect 3180 13626 3236 13628
rect 3260 13626 3316 13628
rect 3340 13626 3396 13628
rect 3420 13626 3476 13628
rect 3180 13574 3226 13626
rect 3226 13574 3236 13626
rect 3260 13574 3290 13626
rect 3290 13574 3302 13626
rect 3302 13574 3316 13626
rect 3340 13574 3354 13626
rect 3354 13574 3366 13626
rect 3366 13574 3396 13626
rect 3420 13574 3430 13626
rect 3430 13574 3476 13626
rect 3180 13572 3236 13574
rect 3260 13572 3316 13574
rect 3340 13572 3396 13574
rect 3420 13572 3476 13574
rect 3180 12538 3236 12540
rect 3260 12538 3316 12540
rect 3340 12538 3396 12540
rect 3420 12538 3476 12540
rect 3180 12486 3226 12538
rect 3226 12486 3236 12538
rect 3260 12486 3290 12538
rect 3290 12486 3302 12538
rect 3302 12486 3316 12538
rect 3340 12486 3354 12538
rect 3354 12486 3366 12538
rect 3366 12486 3396 12538
rect 3420 12486 3430 12538
rect 3430 12486 3476 12538
rect 3180 12484 3236 12486
rect 3260 12484 3316 12486
rect 3340 12484 3396 12486
rect 3420 12484 3476 12486
rect 5404 16346 5460 16348
rect 5484 16346 5540 16348
rect 5564 16346 5620 16348
rect 5644 16346 5700 16348
rect 5404 16294 5450 16346
rect 5450 16294 5460 16346
rect 5484 16294 5514 16346
rect 5514 16294 5526 16346
rect 5526 16294 5540 16346
rect 5564 16294 5578 16346
rect 5578 16294 5590 16346
rect 5590 16294 5620 16346
rect 5644 16294 5654 16346
rect 5654 16294 5700 16346
rect 5404 16292 5460 16294
rect 5484 16292 5540 16294
rect 5564 16292 5620 16294
rect 5644 16292 5700 16294
rect 9852 16346 9908 16348
rect 9932 16346 9988 16348
rect 10012 16346 10068 16348
rect 10092 16346 10148 16348
rect 9852 16294 9898 16346
rect 9898 16294 9908 16346
rect 9932 16294 9962 16346
rect 9962 16294 9974 16346
rect 9974 16294 9988 16346
rect 10012 16294 10026 16346
rect 10026 16294 10038 16346
rect 10038 16294 10068 16346
rect 10092 16294 10102 16346
rect 10102 16294 10148 16346
rect 9852 16292 9908 16294
rect 9932 16292 9988 16294
rect 10012 16292 10068 16294
rect 10092 16292 10148 16294
rect 7628 15802 7684 15804
rect 7708 15802 7764 15804
rect 7788 15802 7844 15804
rect 7868 15802 7924 15804
rect 7628 15750 7674 15802
rect 7674 15750 7684 15802
rect 7708 15750 7738 15802
rect 7738 15750 7750 15802
rect 7750 15750 7764 15802
rect 7788 15750 7802 15802
rect 7802 15750 7814 15802
rect 7814 15750 7844 15802
rect 7868 15750 7878 15802
rect 7878 15750 7924 15802
rect 7628 15748 7684 15750
rect 7708 15748 7764 15750
rect 7788 15748 7844 15750
rect 7868 15748 7924 15750
rect 5404 15258 5460 15260
rect 5484 15258 5540 15260
rect 5564 15258 5620 15260
rect 5644 15258 5700 15260
rect 5404 15206 5450 15258
rect 5450 15206 5460 15258
rect 5484 15206 5514 15258
rect 5514 15206 5526 15258
rect 5526 15206 5540 15258
rect 5564 15206 5578 15258
rect 5578 15206 5590 15258
rect 5590 15206 5620 15258
rect 5644 15206 5654 15258
rect 5654 15206 5700 15258
rect 5404 15204 5460 15206
rect 5484 15204 5540 15206
rect 5564 15204 5620 15206
rect 5644 15204 5700 15206
rect 9852 15258 9908 15260
rect 9932 15258 9988 15260
rect 10012 15258 10068 15260
rect 10092 15258 10148 15260
rect 9852 15206 9898 15258
rect 9898 15206 9908 15258
rect 9932 15206 9962 15258
rect 9962 15206 9974 15258
rect 9974 15206 9988 15258
rect 10012 15206 10026 15258
rect 10026 15206 10038 15258
rect 10038 15206 10068 15258
rect 10092 15206 10102 15258
rect 10102 15206 10148 15258
rect 9852 15204 9908 15206
rect 9932 15204 9988 15206
rect 10012 15204 10068 15206
rect 10092 15204 10148 15206
rect 7628 14714 7684 14716
rect 7708 14714 7764 14716
rect 7788 14714 7844 14716
rect 7868 14714 7924 14716
rect 7628 14662 7674 14714
rect 7674 14662 7684 14714
rect 7708 14662 7738 14714
rect 7738 14662 7750 14714
rect 7750 14662 7764 14714
rect 7788 14662 7802 14714
rect 7802 14662 7814 14714
rect 7814 14662 7844 14714
rect 7868 14662 7878 14714
rect 7878 14662 7924 14714
rect 7628 14660 7684 14662
rect 7708 14660 7764 14662
rect 7788 14660 7844 14662
rect 7868 14660 7924 14662
rect 5404 14170 5460 14172
rect 5484 14170 5540 14172
rect 5564 14170 5620 14172
rect 5644 14170 5700 14172
rect 5404 14118 5450 14170
rect 5450 14118 5460 14170
rect 5484 14118 5514 14170
rect 5514 14118 5526 14170
rect 5526 14118 5540 14170
rect 5564 14118 5578 14170
rect 5578 14118 5590 14170
rect 5590 14118 5620 14170
rect 5644 14118 5654 14170
rect 5654 14118 5700 14170
rect 5404 14116 5460 14118
rect 5484 14116 5540 14118
rect 5564 14116 5620 14118
rect 5644 14116 5700 14118
rect 9852 14170 9908 14172
rect 9932 14170 9988 14172
rect 10012 14170 10068 14172
rect 10092 14170 10148 14172
rect 9852 14118 9898 14170
rect 9898 14118 9908 14170
rect 9932 14118 9962 14170
rect 9962 14118 9974 14170
rect 9974 14118 9988 14170
rect 10012 14118 10026 14170
rect 10026 14118 10038 14170
rect 10038 14118 10068 14170
rect 10092 14118 10102 14170
rect 10102 14118 10148 14170
rect 9852 14116 9908 14118
rect 9932 14116 9988 14118
rect 10012 14116 10068 14118
rect 10092 14116 10148 14118
rect 7628 13626 7684 13628
rect 7708 13626 7764 13628
rect 7788 13626 7844 13628
rect 7868 13626 7924 13628
rect 7628 13574 7674 13626
rect 7674 13574 7684 13626
rect 7708 13574 7738 13626
rect 7738 13574 7750 13626
rect 7750 13574 7764 13626
rect 7788 13574 7802 13626
rect 7802 13574 7814 13626
rect 7814 13574 7844 13626
rect 7868 13574 7878 13626
rect 7878 13574 7924 13626
rect 7628 13572 7684 13574
rect 7708 13572 7764 13574
rect 7788 13572 7844 13574
rect 7868 13572 7924 13574
rect 5404 13082 5460 13084
rect 5484 13082 5540 13084
rect 5564 13082 5620 13084
rect 5644 13082 5700 13084
rect 5404 13030 5450 13082
rect 5450 13030 5460 13082
rect 5484 13030 5514 13082
rect 5514 13030 5526 13082
rect 5526 13030 5540 13082
rect 5564 13030 5578 13082
rect 5578 13030 5590 13082
rect 5590 13030 5620 13082
rect 5644 13030 5654 13082
rect 5654 13030 5700 13082
rect 5404 13028 5460 13030
rect 5484 13028 5540 13030
rect 5564 13028 5620 13030
rect 5644 13028 5700 13030
rect 9852 13082 9908 13084
rect 9932 13082 9988 13084
rect 10012 13082 10068 13084
rect 10092 13082 10148 13084
rect 9852 13030 9898 13082
rect 9898 13030 9908 13082
rect 9932 13030 9962 13082
rect 9962 13030 9974 13082
rect 9974 13030 9988 13082
rect 10012 13030 10026 13082
rect 10026 13030 10038 13082
rect 10038 13030 10068 13082
rect 10092 13030 10102 13082
rect 10102 13030 10148 13082
rect 9852 13028 9908 13030
rect 9932 13028 9988 13030
rect 10012 13028 10068 13030
rect 10092 13028 10148 13030
rect 7628 12538 7684 12540
rect 7708 12538 7764 12540
rect 7788 12538 7844 12540
rect 7868 12538 7924 12540
rect 7628 12486 7674 12538
rect 7674 12486 7684 12538
rect 7708 12486 7738 12538
rect 7738 12486 7750 12538
rect 7750 12486 7764 12538
rect 7788 12486 7802 12538
rect 7802 12486 7814 12538
rect 7814 12486 7844 12538
rect 7868 12486 7878 12538
rect 7878 12486 7924 12538
rect 7628 12484 7684 12486
rect 7708 12484 7764 12486
rect 7788 12484 7844 12486
rect 7868 12484 7924 12486
rect 5404 11994 5460 11996
rect 5484 11994 5540 11996
rect 5564 11994 5620 11996
rect 5644 11994 5700 11996
rect 5404 11942 5450 11994
rect 5450 11942 5460 11994
rect 5484 11942 5514 11994
rect 5514 11942 5526 11994
rect 5526 11942 5540 11994
rect 5564 11942 5578 11994
rect 5578 11942 5590 11994
rect 5590 11942 5620 11994
rect 5644 11942 5654 11994
rect 5654 11942 5700 11994
rect 5404 11940 5460 11942
rect 5484 11940 5540 11942
rect 5564 11940 5620 11942
rect 5644 11940 5700 11942
rect 9852 11994 9908 11996
rect 9932 11994 9988 11996
rect 10012 11994 10068 11996
rect 10092 11994 10148 11996
rect 9852 11942 9898 11994
rect 9898 11942 9908 11994
rect 9932 11942 9962 11994
rect 9962 11942 9974 11994
rect 9974 11942 9988 11994
rect 10012 11942 10026 11994
rect 10026 11942 10038 11994
rect 10038 11942 10068 11994
rect 10092 11942 10102 11994
rect 10102 11942 10148 11994
rect 9852 11940 9908 11942
rect 9932 11940 9988 11942
rect 10012 11940 10068 11942
rect 10092 11940 10148 11942
rect 12076 16890 12132 16892
rect 12156 16890 12212 16892
rect 12236 16890 12292 16892
rect 12316 16890 12372 16892
rect 12076 16838 12122 16890
rect 12122 16838 12132 16890
rect 12156 16838 12186 16890
rect 12186 16838 12198 16890
rect 12198 16838 12212 16890
rect 12236 16838 12250 16890
rect 12250 16838 12262 16890
rect 12262 16838 12292 16890
rect 12316 16838 12326 16890
rect 12326 16838 12372 16890
rect 12076 16836 12132 16838
rect 12156 16836 12212 16838
rect 12236 16836 12292 16838
rect 12316 16836 12372 16838
rect 16524 16890 16580 16892
rect 16604 16890 16660 16892
rect 16684 16890 16740 16892
rect 16764 16890 16820 16892
rect 16524 16838 16570 16890
rect 16570 16838 16580 16890
rect 16604 16838 16634 16890
rect 16634 16838 16646 16890
rect 16646 16838 16660 16890
rect 16684 16838 16698 16890
rect 16698 16838 16710 16890
rect 16710 16838 16740 16890
rect 16764 16838 16774 16890
rect 16774 16838 16820 16890
rect 16524 16836 16580 16838
rect 16604 16836 16660 16838
rect 16684 16836 16740 16838
rect 16764 16836 16820 16838
rect 14300 16346 14356 16348
rect 14380 16346 14436 16348
rect 14460 16346 14516 16348
rect 14540 16346 14596 16348
rect 14300 16294 14346 16346
rect 14346 16294 14356 16346
rect 14380 16294 14410 16346
rect 14410 16294 14422 16346
rect 14422 16294 14436 16346
rect 14460 16294 14474 16346
rect 14474 16294 14486 16346
rect 14486 16294 14516 16346
rect 14540 16294 14550 16346
rect 14550 16294 14596 16346
rect 14300 16292 14356 16294
rect 14380 16292 14436 16294
rect 14460 16292 14516 16294
rect 14540 16292 14596 16294
rect 12076 15802 12132 15804
rect 12156 15802 12212 15804
rect 12236 15802 12292 15804
rect 12316 15802 12372 15804
rect 12076 15750 12122 15802
rect 12122 15750 12132 15802
rect 12156 15750 12186 15802
rect 12186 15750 12198 15802
rect 12198 15750 12212 15802
rect 12236 15750 12250 15802
rect 12250 15750 12262 15802
rect 12262 15750 12292 15802
rect 12316 15750 12326 15802
rect 12326 15750 12372 15802
rect 12076 15748 12132 15750
rect 12156 15748 12212 15750
rect 12236 15748 12292 15750
rect 12316 15748 12372 15750
rect 16524 15802 16580 15804
rect 16604 15802 16660 15804
rect 16684 15802 16740 15804
rect 16764 15802 16820 15804
rect 16524 15750 16570 15802
rect 16570 15750 16580 15802
rect 16604 15750 16634 15802
rect 16634 15750 16646 15802
rect 16646 15750 16660 15802
rect 16684 15750 16698 15802
rect 16698 15750 16710 15802
rect 16710 15750 16740 15802
rect 16764 15750 16774 15802
rect 16774 15750 16820 15802
rect 16524 15748 16580 15750
rect 16604 15748 16660 15750
rect 16684 15748 16740 15750
rect 16764 15748 16820 15750
rect 14300 15258 14356 15260
rect 14380 15258 14436 15260
rect 14460 15258 14516 15260
rect 14540 15258 14596 15260
rect 14300 15206 14346 15258
rect 14346 15206 14356 15258
rect 14380 15206 14410 15258
rect 14410 15206 14422 15258
rect 14422 15206 14436 15258
rect 14460 15206 14474 15258
rect 14474 15206 14486 15258
rect 14486 15206 14516 15258
rect 14540 15206 14550 15258
rect 14550 15206 14596 15258
rect 14300 15204 14356 15206
rect 14380 15204 14436 15206
rect 14460 15204 14516 15206
rect 14540 15204 14596 15206
rect 12076 14714 12132 14716
rect 12156 14714 12212 14716
rect 12236 14714 12292 14716
rect 12316 14714 12372 14716
rect 12076 14662 12122 14714
rect 12122 14662 12132 14714
rect 12156 14662 12186 14714
rect 12186 14662 12198 14714
rect 12198 14662 12212 14714
rect 12236 14662 12250 14714
rect 12250 14662 12262 14714
rect 12262 14662 12292 14714
rect 12316 14662 12326 14714
rect 12326 14662 12372 14714
rect 12076 14660 12132 14662
rect 12156 14660 12212 14662
rect 12236 14660 12292 14662
rect 12316 14660 12372 14662
rect 16524 14714 16580 14716
rect 16604 14714 16660 14716
rect 16684 14714 16740 14716
rect 16764 14714 16820 14716
rect 16524 14662 16570 14714
rect 16570 14662 16580 14714
rect 16604 14662 16634 14714
rect 16634 14662 16646 14714
rect 16646 14662 16660 14714
rect 16684 14662 16698 14714
rect 16698 14662 16710 14714
rect 16710 14662 16740 14714
rect 16764 14662 16774 14714
rect 16774 14662 16820 14714
rect 16524 14660 16580 14662
rect 16604 14660 16660 14662
rect 16684 14660 16740 14662
rect 16764 14660 16820 14662
rect 14300 14170 14356 14172
rect 14380 14170 14436 14172
rect 14460 14170 14516 14172
rect 14540 14170 14596 14172
rect 14300 14118 14346 14170
rect 14346 14118 14356 14170
rect 14380 14118 14410 14170
rect 14410 14118 14422 14170
rect 14422 14118 14436 14170
rect 14460 14118 14474 14170
rect 14474 14118 14486 14170
rect 14486 14118 14516 14170
rect 14540 14118 14550 14170
rect 14550 14118 14596 14170
rect 14300 14116 14356 14118
rect 14380 14116 14436 14118
rect 14460 14116 14516 14118
rect 14540 14116 14596 14118
rect 12076 13626 12132 13628
rect 12156 13626 12212 13628
rect 12236 13626 12292 13628
rect 12316 13626 12372 13628
rect 12076 13574 12122 13626
rect 12122 13574 12132 13626
rect 12156 13574 12186 13626
rect 12186 13574 12198 13626
rect 12198 13574 12212 13626
rect 12236 13574 12250 13626
rect 12250 13574 12262 13626
rect 12262 13574 12292 13626
rect 12316 13574 12326 13626
rect 12326 13574 12372 13626
rect 12076 13572 12132 13574
rect 12156 13572 12212 13574
rect 12236 13572 12292 13574
rect 12316 13572 12372 13574
rect 16524 13626 16580 13628
rect 16604 13626 16660 13628
rect 16684 13626 16740 13628
rect 16764 13626 16820 13628
rect 16524 13574 16570 13626
rect 16570 13574 16580 13626
rect 16604 13574 16634 13626
rect 16634 13574 16646 13626
rect 16646 13574 16660 13626
rect 16684 13574 16698 13626
rect 16698 13574 16710 13626
rect 16710 13574 16740 13626
rect 16764 13574 16774 13626
rect 16774 13574 16820 13626
rect 16524 13572 16580 13574
rect 16604 13572 16660 13574
rect 16684 13572 16740 13574
rect 16764 13572 16820 13574
rect 14300 13082 14356 13084
rect 14380 13082 14436 13084
rect 14460 13082 14516 13084
rect 14540 13082 14596 13084
rect 14300 13030 14346 13082
rect 14346 13030 14356 13082
rect 14380 13030 14410 13082
rect 14410 13030 14422 13082
rect 14422 13030 14436 13082
rect 14460 13030 14474 13082
rect 14474 13030 14486 13082
rect 14486 13030 14516 13082
rect 14540 13030 14550 13082
rect 14550 13030 14596 13082
rect 14300 13028 14356 13030
rect 14380 13028 14436 13030
rect 14460 13028 14516 13030
rect 14540 13028 14596 13030
rect 12076 12538 12132 12540
rect 12156 12538 12212 12540
rect 12236 12538 12292 12540
rect 12316 12538 12372 12540
rect 12076 12486 12122 12538
rect 12122 12486 12132 12538
rect 12156 12486 12186 12538
rect 12186 12486 12198 12538
rect 12198 12486 12212 12538
rect 12236 12486 12250 12538
rect 12250 12486 12262 12538
rect 12262 12486 12292 12538
rect 12316 12486 12326 12538
rect 12326 12486 12372 12538
rect 12076 12484 12132 12486
rect 12156 12484 12212 12486
rect 12236 12484 12292 12486
rect 12316 12484 12372 12486
rect 16524 12538 16580 12540
rect 16604 12538 16660 12540
rect 16684 12538 16740 12540
rect 16764 12538 16820 12540
rect 16524 12486 16570 12538
rect 16570 12486 16580 12538
rect 16604 12486 16634 12538
rect 16634 12486 16646 12538
rect 16646 12486 16660 12538
rect 16684 12486 16698 12538
rect 16698 12486 16710 12538
rect 16710 12486 16740 12538
rect 16764 12486 16774 12538
rect 16774 12486 16820 12538
rect 16524 12484 16580 12486
rect 16604 12484 16660 12486
rect 16684 12484 16740 12486
rect 16764 12484 16820 12486
rect 3180 11450 3236 11452
rect 3260 11450 3316 11452
rect 3340 11450 3396 11452
rect 3420 11450 3476 11452
rect 3180 11398 3226 11450
rect 3226 11398 3236 11450
rect 3260 11398 3290 11450
rect 3290 11398 3302 11450
rect 3302 11398 3316 11450
rect 3340 11398 3354 11450
rect 3354 11398 3366 11450
rect 3366 11398 3396 11450
rect 3420 11398 3430 11450
rect 3430 11398 3476 11450
rect 3180 11396 3236 11398
rect 3260 11396 3316 11398
rect 3340 11396 3396 11398
rect 3420 11396 3476 11398
rect 7628 11450 7684 11452
rect 7708 11450 7764 11452
rect 7788 11450 7844 11452
rect 7868 11450 7924 11452
rect 7628 11398 7674 11450
rect 7674 11398 7684 11450
rect 7708 11398 7738 11450
rect 7738 11398 7750 11450
rect 7750 11398 7764 11450
rect 7788 11398 7802 11450
rect 7802 11398 7814 11450
rect 7814 11398 7844 11450
rect 7868 11398 7878 11450
rect 7878 11398 7924 11450
rect 7628 11396 7684 11398
rect 7708 11396 7764 11398
rect 7788 11396 7844 11398
rect 7868 11396 7924 11398
rect 5404 10906 5460 10908
rect 5484 10906 5540 10908
rect 5564 10906 5620 10908
rect 5644 10906 5700 10908
rect 5404 10854 5450 10906
rect 5450 10854 5460 10906
rect 5484 10854 5514 10906
rect 5514 10854 5526 10906
rect 5526 10854 5540 10906
rect 5564 10854 5578 10906
rect 5578 10854 5590 10906
rect 5590 10854 5620 10906
rect 5644 10854 5654 10906
rect 5654 10854 5700 10906
rect 5404 10852 5460 10854
rect 5484 10852 5540 10854
rect 5564 10852 5620 10854
rect 5644 10852 5700 10854
rect 9852 10906 9908 10908
rect 9932 10906 9988 10908
rect 10012 10906 10068 10908
rect 10092 10906 10148 10908
rect 9852 10854 9898 10906
rect 9898 10854 9908 10906
rect 9932 10854 9962 10906
rect 9962 10854 9974 10906
rect 9974 10854 9988 10906
rect 10012 10854 10026 10906
rect 10026 10854 10038 10906
rect 10038 10854 10068 10906
rect 10092 10854 10102 10906
rect 10102 10854 10148 10906
rect 9852 10852 9908 10854
rect 9932 10852 9988 10854
rect 10012 10852 10068 10854
rect 10092 10852 10148 10854
rect 3180 10362 3236 10364
rect 3260 10362 3316 10364
rect 3340 10362 3396 10364
rect 3420 10362 3476 10364
rect 3180 10310 3226 10362
rect 3226 10310 3236 10362
rect 3260 10310 3290 10362
rect 3290 10310 3302 10362
rect 3302 10310 3316 10362
rect 3340 10310 3354 10362
rect 3354 10310 3366 10362
rect 3366 10310 3396 10362
rect 3420 10310 3430 10362
rect 3430 10310 3476 10362
rect 3180 10308 3236 10310
rect 3260 10308 3316 10310
rect 3340 10308 3396 10310
rect 3420 10308 3476 10310
rect 7628 10362 7684 10364
rect 7708 10362 7764 10364
rect 7788 10362 7844 10364
rect 7868 10362 7924 10364
rect 7628 10310 7674 10362
rect 7674 10310 7684 10362
rect 7708 10310 7738 10362
rect 7738 10310 7750 10362
rect 7750 10310 7764 10362
rect 7788 10310 7802 10362
rect 7802 10310 7814 10362
rect 7814 10310 7844 10362
rect 7868 10310 7878 10362
rect 7878 10310 7924 10362
rect 7628 10308 7684 10310
rect 7708 10308 7764 10310
rect 7788 10308 7844 10310
rect 7868 10308 7924 10310
rect 5404 9818 5460 9820
rect 5484 9818 5540 9820
rect 5564 9818 5620 9820
rect 5644 9818 5700 9820
rect 5404 9766 5450 9818
rect 5450 9766 5460 9818
rect 5484 9766 5514 9818
rect 5514 9766 5526 9818
rect 5526 9766 5540 9818
rect 5564 9766 5578 9818
rect 5578 9766 5590 9818
rect 5590 9766 5620 9818
rect 5644 9766 5654 9818
rect 5654 9766 5700 9818
rect 5404 9764 5460 9766
rect 5484 9764 5540 9766
rect 5564 9764 5620 9766
rect 5644 9764 5700 9766
rect 9852 9818 9908 9820
rect 9932 9818 9988 9820
rect 10012 9818 10068 9820
rect 10092 9818 10148 9820
rect 9852 9766 9898 9818
rect 9898 9766 9908 9818
rect 9932 9766 9962 9818
rect 9962 9766 9974 9818
rect 9974 9766 9988 9818
rect 10012 9766 10026 9818
rect 10026 9766 10038 9818
rect 10038 9766 10068 9818
rect 10092 9766 10102 9818
rect 10102 9766 10148 9818
rect 9852 9764 9908 9766
rect 9932 9764 9988 9766
rect 10012 9764 10068 9766
rect 10092 9764 10148 9766
rect 3180 9274 3236 9276
rect 3260 9274 3316 9276
rect 3340 9274 3396 9276
rect 3420 9274 3476 9276
rect 3180 9222 3226 9274
rect 3226 9222 3236 9274
rect 3260 9222 3290 9274
rect 3290 9222 3302 9274
rect 3302 9222 3316 9274
rect 3340 9222 3354 9274
rect 3354 9222 3366 9274
rect 3366 9222 3396 9274
rect 3420 9222 3430 9274
rect 3430 9222 3476 9274
rect 3180 9220 3236 9222
rect 3260 9220 3316 9222
rect 3340 9220 3396 9222
rect 3420 9220 3476 9222
rect 7628 9274 7684 9276
rect 7708 9274 7764 9276
rect 7788 9274 7844 9276
rect 7868 9274 7924 9276
rect 7628 9222 7674 9274
rect 7674 9222 7684 9274
rect 7708 9222 7738 9274
rect 7738 9222 7750 9274
rect 7750 9222 7764 9274
rect 7788 9222 7802 9274
rect 7802 9222 7814 9274
rect 7814 9222 7844 9274
rect 7868 9222 7878 9274
rect 7878 9222 7924 9274
rect 7628 9220 7684 9222
rect 7708 9220 7764 9222
rect 7788 9220 7844 9222
rect 7868 9220 7924 9222
rect 5404 8730 5460 8732
rect 5484 8730 5540 8732
rect 5564 8730 5620 8732
rect 5644 8730 5700 8732
rect 5404 8678 5450 8730
rect 5450 8678 5460 8730
rect 5484 8678 5514 8730
rect 5514 8678 5526 8730
rect 5526 8678 5540 8730
rect 5564 8678 5578 8730
rect 5578 8678 5590 8730
rect 5590 8678 5620 8730
rect 5644 8678 5654 8730
rect 5654 8678 5700 8730
rect 5404 8676 5460 8678
rect 5484 8676 5540 8678
rect 5564 8676 5620 8678
rect 5644 8676 5700 8678
rect 9852 8730 9908 8732
rect 9932 8730 9988 8732
rect 10012 8730 10068 8732
rect 10092 8730 10148 8732
rect 9852 8678 9898 8730
rect 9898 8678 9908 8730
rect 9932 8678 9962 8730
rect 9962 8678 9974 8730
rect 9974 8678 9988 8730
rect 10012 8678 10026 8730
rect 10026 8678 10038 8730
rect 10038 8678 10068 8730
rect 10092 8678 10102 8730
rect 10102 8678 10148 8730
rect 9852 8676 9908 8678
rect 9932 8676 9988 8678
rect 10012 8676 10068 8678
rect 10092 8676 10148 8678
rect 3180 8186 3236 8188
rect 3260 8186 3316 8188
rect 3340 8186 3396 8188
rect 3420 8186 3476 8188
rect 3180 8134 3226 8186
rect 3226 8134 3236 8186
rect 3260 8134 3290 8186
rect 3290 8134 3302 8186
rect 3302 8134 3316 8186
rect 3340 8134 3354 8186
rect 3354 8134 3366 8186
rect 3366 8134 3396 8186
rect 3420 8134 3430 8186
rect 3430 8134 3476 8186
rect 3180 8132 3236 8134
rect 3260 8132 3316 8134
rect 3340 8132 3396 8134
rect 3420 8132 3476 8134
rect 7628 8186 7684 8188
rect 7708 8186 7764 8188
rect 7788 8186 7844 8188
rect 7868 8186 7924 8188
rect 7628 8134 7674 8186
rect 7674 8134 7684 8186
rect 7708 8134 7738 8186
rect 7738 8134 7750 8186
rect 7750 8134 7764 8186
rect 7788 8134 7802 8186
rect 7802 8134 7814 8186
rect 7814 8134 7844 8186
rect 7868 8134 7878 8186
rect 7878 8134 7924 8186
rect 7628 8132 7684 8134
rect 7708 8132 7764 8134
rect 7788 8132 7844 8134
rect 7868 8132 7924 8134
rect 14300 11994 14356 11996
rect 14380 11994 14436 11996
rect 14460 11994 14516 11996
rect 14540 11994 14596 11996
rect 14300 11942 14346 11994
rect 14346 11942 14356 11994
rect 14380 11942 14410 11994
rect 14410 11942 14422 11994
rect 14422 11942 14436 11994
rect 14460 11942 14474 11994
rect 14474 11942 14486 11994
rect 14486 11942 14516 11994
rect 14540 11942 14550 11994
rect 14550 11942 14596 11994
rect 14300 11940 14356 11942
rect 14380 11940 14436 11942
rect 14460 11940 14516 11942
rect 14540 11940 14596 11942
rect 12076 11450 12132 11452
rect 12156 11450 12212 11452
rect 12236 11450 12292 11452
rect 12316 11450 12372 11452
rect 12076 11398 12122 11450
rect 12122 11398 12132 11450
rect 12156 11398 12186 11450
rect 12186 11398 12198 11450
rect 12198 11398 12212 11450
rect 12236 11398 12250 11450
rect 12250 11398 12262 11450
rect 12262 11398 12292 11450
rect 12316 11398 12326 11450
rect 12326 11398 12372 11450
rect 12076 11396 12132 11398
rect 12156 11396 12212 11398
rect 12236 11396 12292 11398
rect 12316 11396 12372 11398
rect 12076 10362 12132 10364
rect 12156 10362 12212 10364
rect 12236 10362 12292 10364
rect 12316 10362 12372 10364
rect 12076 10310 12122 10362
rect 12122 10310 12132 10362
rect 12156 10310 12186 10362
rect 12186 10310 12198 10362
rect 12198 10310 12212 10362
rect 12236 10310 12250 10362
rect 12250 10310 12262 10362
rect 12262 10310 12292 10362
rect 12316 10310 12326 10362
rect 12326 10310 12372 10362
rect 12076 10308 12132 10310
rect 12156 10308 12212 10310
rect 12236 10308 12292 10310
rect 12316 10308 12372 10310
rect 18142 11600 18198 11656
rect 16524 11450 16580 11452
rect 16604 11450 16660 11452
rect 16684 11450 16740 11452
rect 16764 11450 16820 11452
rect 16524 11398 16570 11450
rect 16570 11398 16580 11450
rect 16604 11398 16634 11450
rect 16634 11398 16646 11450
rect 16646 11398 16660 11450
rect 16684 11398 16698 11450
rect 16698 11398 16710 11450
rect 16710 11398 16740 11450
rect 16764 11398 16774 11450
rect 16774 11398 16820 11450
rect 16524 11396 16580 11398
rect 16604 11396 16660 11398
rect 16684 11396 16740 11398
rect 16764 11396 16820 11398
rect 14300 10906 14356 10908
rect 14380 10906 14436 10908
rect 14460 10906 14516 10908
rect 14540 10906 14596 10908
rect 14300 10854 14346 10906
rect 14346 10854 14356 10906
rect 14380 10854 14410 10906
rect 14410 10854 14422 10906
rect 14422 10854 14436 10906
rect 14460 10854 14474 10906
rect 14474 10854 14486 10906
rect 14486 10854 14516 10906
rect 14540 10854 14550 10906
rect 14550 10854 14596 10906
rect 14300 10852 14356 10854
rect 14380 10852 14436 10854
rect 14460 10852 14516 10854
rect 14540 10852 14596 10854
rect 14300 9818 14356 9820
rect 14380 9818 14436 9820
rect 14460 9818 14516 9820
rect 14540 9818 14596 9820
rect 14300 9766 14346 9818
rect 14346 9766 14356 9818
rect 14380 9766 14410 9818
rect 14410 9766 14422 9818
rect 14422 9766 14436 9818
rect 14460 9766 14474 9818
rect 14474 9766 14486 9818
rect 14486 9766 14516 9818
rect 14540 9766 14550 9818
rect 14550 9766 14596 9818
rect 14300 9764 14356 9766
rect 14380 9764 14436 9766
rect 14460 9764 14516 9766
rect 14540 9764 14596 9766
rect 12076 9274 12132 9276
rect 12156 9274 12212 9276
rect 12236 9274 12292 9276
rect 12316 9274 12372 9276
rect 12076 9222 12122 9274
rect 12122 9222 12132 9274
rect 12156 9222 12186 9274
rect 12186 9222 12198 9274
rect 12198 9222 12212 9274
rect 12236 9222 12250 9274
rect 12250 9222 12262 9274
rect 12262 9222 12292 9274
rect 12316 9222 12326 9274
rect 12326 9222 12372 9274
rect 12076 9220 12132 9222
rect 12156 9220 12212 9222
rect 12236 9220 12292 9222
rect 12316 9220 12372 9222
rect 14300 8730 14356 8732
rect 14380 8730 14436 8732
rect 14460 8730 14516 8732
rect 14540 8730 14596 8732
rect 14300 8678 14346 8730
rect 14346 8678 14356 8730
rect 14380 8678 14410 8730
rect 14410 8678 14422 8730
rect 14422 8678 14436 8730
rect 14460 8678 14474 8730
rect 14474 8678 14486 8730
rect 14486 8678 14516 8730
rect 14540 8678 14550 8730
rect 14550 8678 14596 8730
rect 14300 8676 14356 8678
rect 14380 8676 14436 8678
rect 14460 8676 14516 8678
rect 14540 8676 14596 8678
rect 12076 8186 12132 8188
rect 12156 8186 12212 8188
rect 12236 8186 12292 8188
rect 12316 8186 12372 8188
rect 12076 8134 12122 8186
rect 12122 8134 12132 8186
rect 12156 8134 12186 8186
rect 12186 8134 12198 8186
rect 12198 8134 12212 8186
rect 12236 8134 12250 8186
rect 12250 8134 12262 8186
rect 12262 8134 12292 8186
rect 12316 8134 12326 8186
rect 12326 8134 12372 8186
rect 12076 8132 12132 8134
rect 12156 8132 12212 8134
rect 12236 8132 12292 8134
rect 12316 8132 12372 8134
rect 5404 7642 5460 7644
rect 5484 7642 5540 7644
rect 5564 7642 5620 7644
rect 5644 7642 5700 7644
rect 5404 7590 5450 7642
rect 5450 7590 5460 7642
rect 5484 7590 5514 7642
rect 5514 7590 5526 7642
rect 5526 7590 5540 7642
rect 5564 7590 5578 7642
rect 5578 7590 5590 7642
rect 5590 7590 5620 7642
rect 5644 7590 5654 7642
rect 5654 7590 5700 7642
rect 5404 7588 5460 7590
rect 5484 7588 5540 7590
rect 5564 7588 5620 7590
rect 5644 7588 5700 7590
rect 9852 7642 9908 7644
rect 9932 7642 9988 7644
rect 10012 7642 10068 7644
rect 10092 7642 10148 7644
rect 9852 7590 9898 7642
rect 9898 7590 9908 7642
rect 9932 7590 9962 7642
rect 9962 7590 9974 7642
rect 9974 7590 9988 7642
rect 10012 7590 10026 7642
rect 10026 7590 10038 7642
rect 10038 7590 10068 7642
rect 10092 7590 10102 7642
rect 10102 7590 10148 7642
rect 9852 7588 9908 7590
rect 9932 7588 9988 7590
rect 10012 7588 10068 7590
rect 10092 7588 10148 7590
rect 14300 7642 14356 7644
rect 14380 7642 14436 7644
rect 14460 7642 14516 7644
rect 14540 7642 14596 7644
rect 14300 7590 14346 7642
rect 14346 7590 14356 7642
rect 14380 7590 14410 7642
rect 14410 7590 14422 7642
rect 14422 7590 14436 7642
rect 14460 7590 14474 7642
rect 14474 7590 14486 7642
rect 14486 7590 14516 7642
rect 14540 7590 14550 7642
rect 14550 7590 14596 7642
rect 14300 7588 14356 7590
rect 14380 7588 14436 7590
rect 14460 7588 14516 7590
rect 14540 7588 14596 7590
rect 3180 7098 3236 7100
rect 3260 7098 3316 7100
rect 3340 7098 3396 7100
rect 3420 7098 3476 7100
rect 3180 7046 3226 7098
rect 3226 7046 3236 7098
rect 3260 7046 3290 7098
rect 3290 7046 3302 7098
rect 3302 7046 3316 7098
rect 3340 7046 3354 7098
rect 3354 7046 3366 7098
rect 3366 7046 3396 7098
rect 3420 7046 3430 7098
rect 3430 7046 3476 7098
rect 3180 7044 3236 7046
rect 3260 7044 3316 7046
rect 3340 7044 3396 7046
rect 3420 7044 3476 7046
rect 7628 7098 7684 7100
rect 7708 7098 7764 7100
rect 7788 7098 7844 7100
rect 7868 7098 7924 7100
rect 7628 7046 7674 7098
rect 7674 7046 7684 7098
rect 7708 7046 7738 7098
rect 7738 7046 7750 7098
rect 7750 7046 7764 7098
rect 7788 7046 7802 7098
rect 7802 7046 7814 7098
rect 7814 7046 7844 7098
rect 7868 7046 7878 7098
rect 7878 7046 7924 7098
rect 7628 7044 7684 7046
rect 7708 7044 7764 7046
rect 7788 7044 7844 7046
rect 7868 7044 7924 7046
rect 12076 7098 12132 7100
rect 12156 7098 12212 7100
rect 12236 7098 12292 7100
rect 12316 7098 12372 7100
rect 12076 7046 12122 7098
rect 12122 7046 12132 7098
rect 12156 7046 12186 7098
rect 12186 7046 12198 7098
rect 12198 7046 12212 7098
rect 12236 7046 12250 7098
rect 12250 7046 12262 7098
rect 12262 7046 12292 7098
rect 12316 7046 12326 7098
rect 12326 7046 12372 7098
rect 12076 7044 12132 7046
rect 12156 7044 12212 7046
rect 12236 7044 12292 7046
rect 12316 7044 12372 7046
rect 5404 6554 5460 6556
rect 5484 6554 5540 6556
rect 5564 6554 5620 6556
rect 5644 6554 5700 6556
rect 5404 6502 5450 6554
rect 5450 6502 5460 6554
rect 5484 6502 5514 6554
rect 5514 6502 5526 6554
rect 5526 6502 5540 6554
rect 5564 6502 5578 6554
rect 5578 6502 5590 6554
rect 5590 6502 5620 6554
rect 5644 6502 5654 6554
rect 5654 6502 5700 6554
rect 5404 6500 5460 6502
rect 5484 6500 5540 6502
rect 5564 6500 5620 6502
rect 5644 6500 5700 6502
rect 9852 6554 9908 6556
rect 9932 6554 9988 6556
rect 10012 6554 10068 6556
rect 10092 6554 10148 6556
rect 9852 6502 9898 6554
rect 9898 6502 9908 6554
rect 9932 6502 9962 6554
rect 9962 6502 9974 6554
rect 9974 6502 9988 6554
rect 10012 6502 10026 6554
rect 10026 6502 10038 6554
rect 10038 6502 10068 6554
rect 10092 6502 10102 6554
rect 10102 6502 10148 6554
rect 9852 6500 9908 6502
rect 9932 6500 9988 6502
rect 10012 6500 10068 6502
rect 10092 6500 10148 6502
rect 14300 6554 14356 6556
rect 14380 6554 14436 6556
rect 14460 6554 14516 6556
rect 14540 6554 14596 6556
rect 14300 6502 14346 6554
rect 14346 6502 14356 6554
rect 14380 6502 14410 6554
rect 14410 6502 14422 6554
rect 14422 6502 14436 6554
rect 14460 6502 14474 6554
rect 14474 6502 14486 6554
rect 14486 6502 14516 6554
rect 14540 6502 14550 6554
rect 14550 6502 14596 6554
rect 14300 6500 14356 6502
rect 14380 6500 14436 6502
rect 14460 6500 14516 6502
rect 14540 6500 14596 6502
rect 3180 6010 3236 6012
rect 3260 6010 3316 6012
rect 3340 6010 3396 6012
rect 3420 6010 3476 6012
rect 3180 5958 3226 6010
rect 3226 5958 3236 6010
rect 3260 5958 3290 6010
rect 3290 5958 3302 6010
rect 3302 5958 3316 6010
rect 3340 5958 3354 6010
rect 3354 5958 3366 6010
rect 3366 5958 3396 6010
rect 3420 5958 3430 6010
rect 3430 5958 3476 6010
rect 3180 5956 3236 5958
rect 3260 5956 3316 5958
rect 3340 5956 3396 5958
rect 3420 5956 3476 5958
rect 7628 6010 7684 6012
rect 7708 6010 7764 6012
rect 7788 6010 7844 6012
rect 7868 6010 7924 6012
rect 7628 5958 7674 6010
rect 7674 5958 7684 6010
rect 7708 5958 7738 6010
rect 7738 5958 7750 6010
rect 7750 5958 7764 6010
rect 7788 5958 7802 6010
rect 7802 5958 7814 6010
rect 7814 5958 7844 6010
rect 7868 5958 7878 6010
rect 7878 5958 7924 6010
rect 7628 5956 7684 5958
rect 7708 5956 7764 5958
rect 7788 5956 7844 5958
rect 7868 5956 7924 5958
rect 12076 6010 12132 6012
rect 12156 6010 12212 6012
rect 12236 6010 12292 6012
rect 12316 6010 12372 6012
rect 12076 5958 12122 6010
rect 12122 5958 12132 6010
rect 12156 5958 12186 6010
rect 12186 5958 12198 6010
rect 12198 5958 12212 6010
rect 12236 5958 12250 6010
rect 12250 5958 12262 6010
rect 12262 5958 12292 6010
rect 12316 5958 12326 6010
rect 12326 5958 12372 6010
rect 12076 5956 12132 5958
rect 12156 5956 12212 5958
rect 12236 5956 12292 5958
rect 12316 5956 12372 5958
rect 5404 5466 5460 5468
rect 5484 5466 5540 5468
rect 5564 5466 5620 5468
rect 5644 5466 5700 5468
rect 5404 5414 5450 5466
rect 5450 5414 5460 5466
rect 5484 5414 5514 5466
rect 5514 5414 5526 5466
rect 5526 5414 5540 5466
rect 5564 5414 5578 5466
rect 5578 5414 5590 5466
rect 5590 5414 5620 5466
rect 5644 5414 5654 5466
rect 5654 5414 5700 5466
rect 5404 5412 5460 5414
rect 5484 5412 5540 5414
rect 5564 5412 5620 5414
rect 5644 5412 5700 5414
rect 9852 5466 9908 5468
rect 9932 5466 9988 5468
rect 10012 5466 10068 5468
rect 10092 5466 10148 5468
rect 9852 5414 9898 5466
rect 9898 5414 9908 5466
rect 9932 5414 9962 5466
rect 9962 5414 9974 5466
rect 9974 5414 9988 5466
rect 10012 5414 10026 5466
rect 10026 5414 10038 5466
rect 10038 5414 10068 5466
rect 10092 5414 10102 5466
rect 10102 5414 10148 5466
rect 9852 5412 9908 5414
rect 9932 5412 9988 5414
rect 10012 5412 10068 5414
rect 10092 5412 10148 5414
rect 14300 5466 14356 5468
rect 14380 5466 14436 5468
rect 14460 5466 14516 5468
rect 14540 5466 14596 5468
rect 14300 5414 14346 5466
rect 14346 5414 14356 5466
rect 14380 5414 14410 5466
rect 14410 5414 14422 5466
rect 14422 5414 14436 5466
rect 14460 5414 14474 5466
rect 14474 5414 14486 5466
rect 14486 5414 14516 5466
rect 14540 5414 14550 5466
rect 14550 5414 14596 5466
rect 14300 5412 14356 5414
rect 14380 5412 14436 5414
rect 14460 5412 14516 5414
rect 14540 5412 14596 5414
rect 3180 4922 3236 4924
rect 3260 4922 3316 4924
rect 3340 4922 3396 4924
rect 3420 4922 3476 4924
rect 3180 4870 3226 4922
rect 3226 4870 3236 4922
rect 3260 4870 3290 4922
rect 3290 4870 3302 4922
rect 3302 4870 3316 4922
rect 3340 4870 3354 4922
rect 3354 4870 3366 4922
rect 3366 4870 3396 4922
rect 3420 4870 3430 4922
rect 3430 4870 3476 4922
rect 3180 4868 3236 4870
rect 3260 4868 3316 4870
rect 3340 4868 3396 4870
rect 3420 4868 3476 4870
rect 7628 4922 7684 4924
rect 7708 4922 7764 4924
rect 7788 4922 7844 4924
rect 7868 4922 7924 4924
rect 7628 4870 7674 4922
rect 7674 4870 7684 4922
rect 7708 4870 7738 4922
rect 7738 4870 7750 4922
rect 7750 4870 7764 4922
rect 7788 4870 7802 4922
rect 7802 4870 7814 4922
rect 7814 4870 7844 4922
rect 7868 4870 7878 4922
rect 7878 4870 7924 4922
rect 7628 4868 7684 4870
rect 7708 4868 7764 4870
rect 7788 4868 7844 4870
rect 7868 4868 7924 4870
rect 12076 4922 12132 4924
rect 12156 4922 12212 4924
rect 12236 4922 12292 4924
rect 12316 4922 12372 4924
rect 12076 4870 12122 4922
rect 12122 4870 12132 4922
rect 12156 4870 12186 4922
rect 12186 4870 12198 4922
rect 12198 4870 12212 4922
rect 12236 4870 12250 4922
rect 12250 4870 12262 4922
rect 12262 4870 12292 4922
rect 12316 4870 12326 4922
rect 12326 4870 12372 4922
rect 12076 4868 12132 4870
rect 12156 4868 12212 4870
rect 12236 4868 12292 4870
rect 12316 4868 12372 4870
rect 5404 4378 5460 4380
rect 5484 4378 5540 4380
rect 5564 4378 5620 4380
rect 5644 4378 5700 4380
rect 5404 4326 5450 4378
rect 5450 4326 5460 4378
rect 5484 4326 5514 4378
rect 5514 4326 5526 4378
rect 5526 4326 5540 4378
rect 5564 4326 5578 4378
rect 5578 4326 5590 4378
rect 5590 4326 5620 4378
rect 5644 4326 5654 4378
rect 5654 4326 5700 4378
rect 5404 4324 5460 4326
rect 5484 4324 5540 4326
rect 5564 4324 5620 4326
rect 5644 4324 5700 4326
rect 9852 4378 9908 4380
rect 9932 4378 9988 4380
rect 10012 4378 10068 4380
rect 10092 4378 10148 4380
rect 9852 4326 9898 4378
rect 9898 4326 9908 4378
rect 9932 4326 9962 4378
rect 9962 4326 9974 4378
rect 9974 4326 9988 4378
rect 10012 4326 10026 4378
rect 10026 4326 10038 4378
rect 10038 4326 10068 4378
rect 10092 4326 10102 4378
rect 10102 4326 10148 4378
rect 9852 4324 9908 4326
rect 9932 4324 9988 4326
rect 10012 4324 10068 4326
rect 10092 4324 10148 4326
rect 14300 4378 14356 4380
rect 14380 4378 14436 4380
rect 14460 4378 14516 4380
rect 14540 4378 14596 4380
rect 14300 4326 14346 4378
rect 14346 4326 14356 4378
rect 14380 4326 14410 4378
rect 14410 4326 14422 4378
rect 14422 4326 14436 4378
rect 14460 4326 14474 4378
rect 14474 4326 14486 4378
rect 14486 4326 14516 4378
rect 14540 4326 14550 4378
rect 14550 4326 14596 4378
rect 14300 4324 14356 4326
rect 14380 4324 14436 4326
rect 14460 4324 14516 4326
rect 14540 4324 14596 4326
rect 3180 3834 3236 3836
rect 3260 3834 3316 3836
rect 3340 3834 3396 3836
rect 3420 3834 3476 3836
rect 3180 3782 3226 3834
rect 3226 3782 3236 3834
rect 3260 3782 3290 3834
rect 3290 3782 3302 3834
rect 3302 3782 3316 3834
rect 3340 3782 3354 3834
rect 3354 3782 3366 3834
rect 3366 3782 3396 3834
rect 3420 3782 3430 3834
rect 3430 3782 3476 3834
rect 3180 3780 3236 3782
rect 3260 3780 3316 3782
rect 3340 3780 3396 3782
rect 3420 3780 3476 3782
rect 7628 3834 7684 3836
rect 7708 3834 7764 3836
rect 7788 3834 7844 3836
rect 7868 3834 7924 3836
rect 7628 3782 7674 3834
rect 7674 3782 7684 3834
rect 7708 3782 7738 3834
rect 7738 3782 7750 3834
rect 7750 3782 7764 3834
rect 7788 3782 7802 3834
rect 7802 3782 7814 3834
rect 7814 3782 7844 3834
rect 7868 3782 7878 3834
rect 7878 3782 7924 3834
rect 7628 3780 7684 3782
rect 7708 3780 7764 3782
rect 7788 3780 7844 3782
rect 7868 3780 7924 3782
rect 12076 3834 12132 3836
rect 12156 3834 12212 3836
rect 12236 3834 12292 3836
rect 12316 3834 12372 3836
rect 12076 3782 12122 3834
rect 12122 3782 12132 3834
rect 12156 3782 12186 3834
rect 12186 3782 12198 3834
rect 12198 3782 12212 3834
rect 12236 3782 12250 3834
rect 12250 3782 12262 3834
rect 12262 3782 12292 3834
rect 12316 3782 12326 3834
rect 12326 3782 12372 3834
rect 12076 3780 12132 3782
rect 12156 3780 12212 3782
rect 12236 3780 12292 3782
rect 12316 3780 12372 3782
rect 5404 3290 5460 3292
rect 5484 3290 5540 3292
rect 5564 3290 5620 3292
rect 5644 3290 5700 3292
rect 5404 3238 5450 3290
rect 5450 3238 5460 3290
rect 5484 3238 5514 3290
rect 5514 3238 5526 3290
rect 5526 3238 5540 3290
rect 5564 3238 5578 3290
rect 5578 3238 5590 3290
rect 5590 3238 5620 3290
rect 5644 3238 5654 3290
rect 5654 3238 5700 3290
rect 5404 3236 5460 3238
rect 5484 3236 5540 3238
rect 5564 3236 5620 3238
rect 5644 3236 5700 3238
rect 9852 3290 9908 3292
rect 9932 3290 9988 3292
rect 10012 3290 10068 3292
rect 10092 3290 10148 3292
rect 9852 3238 9898 3290
rect 9898 3238 9908 3290
rect 9932 3238 9962 3290
rect 9962 3238 9974 3290
rect 9974 3238 9988 3290
rect 10012 3238 10026 3290
rect 10026 3238 10038 3290
rect 10038 3238 10068 3290
rect 10092 3238 10102 3290
rect 10102 3238 10148 3290
rect 9852 3236 9908 3238
rect 9932 3236 9988 3238
rect 10012 3236 10068 3238
rect 10092 3236 10148 3238
rect 14300 3290 14356 3292
rect 14380 3290 14436 3292
rect 14460 3290 14516 3292
rect 14540 3290 14596 3292
rect 14300 3238 14346 3290
rect 14346 3238 14356 3290
rect 14380 3238 14410 3290
rect 14410 3238 14422 3290
rect 14422 3238 14436 3290
rect 14460 3238 14474 3290
rect 14474 3238 14486 3290
rect 14486 3238 14516 3290
rect 14540 3238 14550 3290
rect 14550 3238 14596 3290
rect 14300 3236 14356 3238
rect 14380 3236 14436 3238
rect 14460 3236 14516 3238
rect 14540 3236 14596 3238
rect 3180 2746 3236 2748
rect 3260 2746 3316 2748
rect 3340 2746 3396 2748
rect 3420 2746 3476 2748
rect 3180 2694 3226 2746
rect 3226 2694 3236 2746
rect 3260 2694 3290 2746
rect 3290 2694 3302 2746
rect 3302 2694 3316 2746
rect 3340 2694 3354 2746
rect 3354 2694 3366 2746
rect 3366 2694 3396 2746
rect 3420 2694 3430 2746
rect 3430 2694 3476 2746
rect 3180 2692 3236 2694
rect 3260 2692 3316 2694
rect 3340 2692 3396 2694
rect 3420 2692 3476 2694
rect 7628 2746 7684 2748
rect 7708 2746 7764 2748
rect 7788 2746 7844 2748
rect 7868 2746 7924 2748
rect 7628 2694 7674 2746
rect 7674 2694 7684 2746
rect 7708 2694 7738 2746
rect 7738 2694 7750 2746
rect 7750 2694 7764 2746
rect 7788 2694 7802 2746
rect 7802 2694 7814 2746
rect 7814 2694 7844 2746
rect 7868 2694 7878 2746
rect 7878 2694 7924 2746
rect 7628 2692 7684 2694
rect 7708 2692 7764 2694
rect 7788 2692 7844 2694
rect 7868 2692 7924 2694
rect 12076 2746 12132 2748
rect 12156 2746 12212 2748
rect 12236 2746 12292 2748
rect 12316 2746 12372 2748
rect 12076 2694 12122 2746
rect 12122 2694 12132 2746
rect 12156 2694 12186 2746
rect 12186 2694 12198 2746
rect 12198 2694 12212 2746
rect 12236 2694 12250 2746
rect 12250 2694 12262 2746
rect 12262 2694 12292 2746
rect 12316 2694 12326 2746
rect 12326 2694 12372 2746
rect 12076 2692 12132 2694
rect 12156 2692 12212 2694
rect 12236 2692 12292 2694
rect 12316 2692 12372 2694
rect 16524 10362 16580 10364
rect 16604 10362 16660 10364
rect 16684 10362 16740 10364
rect 16764 10362 16820 10364
rect 16524 10310 16570 10362
rect 16570 10310 16580 10362
rect 16604 10310 16634 10362
rect 16634 10310 16646 10362
rect 16646 10310 16660 10362
rect 16684 10310 16698 10362
rect 16698 10310 16710 10362
rect 16710 10310 16740 10362
rect 16764 10310 16774 10362
rect 16774 10310 16820 10362
rect 16524 10308 16580 10310
rect 16604 10308 16660 10310
rect 16684 10308 16740 10310
rect 16764 10308 16820 10310
rect 16524 9274 16580 9276
rect 16604 9274 16660 9276
rect 16684 9274 16740 9276
rect 16764 9274 16820 9276
rect 16524 9222 16570 9274
rect 16570 9222 16580 9274
rect 16604 9222 16634 9274
rect 16634 9222 16646 9274
rect 16646 9222 16660 9274
rect 16684 9222 16698 9274
rect 16698 9222 16710 9274
rect 16710 9222 16740 9274
rect 16764 9222 16774 9274
rect 16774 9222 16820 9274
rect 16524 9220 16580 9222
rect 16604 9220 16660 9222
rect 16684 9220 16740 9222
rect 16764 9220 16820 9222
rect 16524 8186 16580 8188
rect 16604 8186 16660 8188
rect 16684 8186 16740 8188
rect 16764 8186 16820 8188
rect 16524 8134 16570 8186
rect 16570 8134 16580 8186
rect 16604 8134 16634 8186
rect 16634 8134 16646 8186
rect 16646 8134 16660 8186
rect 16684 8134 16698 8186
rect 16698 8134 16710 8186
rect 16710 8134 16740 8186
rect 16764 8134 16774 8186
rect 16774 8134 16820 8186
rect 16524 8132 16580 8134
rect 16604 8132 16660 8134
rect 16684 8132 16740 8134
rect 16764 8132 16820 8134
rect 16524 7098 16580 7100
rect 16604 7098 16660 7100
rect 16684 7098 16740 7100
rect 16764 7098 16820 7100
rect 16524 7046 16570 7098
rect 16570 7046 16580 7098
rect 16604 7046 16634 7098
rect 16634 7046 16646 7098
rect 16646 7046 16660 7098
rect 16684 7046 16698 7098
rect 16698 7046 16710 7098
rect 16710 7046 16740 7098
rect 16764 7046 16774 7098
rect 16774 7046 16820 7098
rect 16524 7044 16580 7046
rect 16604 7044 16660 7046
rect 16684 7044 16740 7046
rect 16764 7044 16820 7046
rect 16524 6010 16580 6012
rect 16604 6010 16660 6012
rect 16684 6010 16740 6012
rect 16764 6010 16820 6012
rect 16524 5958 16570 6010
rect 16570 5958 16580 6010
rect 16604 5958 16634 6010
rect 16634 5958 16646 6010
rect 16646 5958 16660 6010
rect 16684 5958 16698 6010
rect 16698 5958 16710 6010
rect 16710 5958 16740 6010
rect 16764 5958 16774 6010
rect 16774 5958 16820 6010
rect 16524 5956 16580 5958
rect 16604 5956 16660 5958
rect 16684 5956 16740 5958
rect 16764 5956 16820 5958
rect 16524 4922 16580 4924
rect 16604 4922 16660 4924
rect 16684 4922 16740 4924
rect 16764 4922 16820 4924
rect 16524 4870 16570 4922
rect 16570 4870 16580 4922
rect 16604 4870 16634 4922
rect 16634 4870 16646 4922
rect 16646 4870 16660 4922
rect 16684 4870 16698 4922
rect 16698 4870 16710 4922
rect 16710 4870 16740 4922
rect 16764 4870 16774 4922
rect 16774 4870 16820 4922
rect 16524 4868 16580 4870
rect 16604 4868 16660 4870
rect 16684 4868 16740 4870
rect 16764 4868 16820 4870
rect 16524 3834 16580 3836
rect 16604 3834 16660 3836
rect 16684 3834 16740 3836
rect 16764 3834 16820 3836
rect 16524 3782 16570 3834
rect 16570 3782 16580 3834
rect 16604 3782 16634 3834
rect 16634 3782 16646 3834
rect 16646 3782 16660 3834
rect 16684 3782 16698 3834
rect 16698 3782 16710 3834
rect 16710 3782 16740 3834
rect 16764 3782 16774 3834
rect 16774 3782 16820 3834
rect 16524 3780 16580 3782
rect 16604 3780 16660 3782
rect 16684 3780 16740 3782
rect 16764 3780 16820 3782
rect 16524 2746 16580 2748
rect 16604 2746 16660 2748
rect 16684 2746 16740 2748
rect 16764 2746 16820 2748
rect 16524 2694 16570 2746
rect 16570 2694 16580 2746
rect 16604 2694 16634 2746
rect 16634 2694 16646 2746
rect 16646 2694 16660 2746
rect 16684 2694 16698 2746
rect 16698 2694 16710 2746
rect 16710 2694 16740 2746
rect 16764 2694 16774 2746
rect 16774 2694 16820 2746
rect 16524 2692 16580 2694
rect 16604 2692 16660 2694
rect 16684 2692 16740 2694
rect 16764 2692 16820 2694
rect 5404 2202 5460 2204
rect 5484 2202 5540 2204
rect 5564 2202 5620 2204
rect 5644 2202 5700 2204
rect 5404 2150 5450 2202
rect 5450 2150 5460 2202
rect 5484 2150 5514 2202
rect 5514 2150 5526 2202
rect 5526 2150 5540 2202
rect 5564 2150 5578 2202
rect 5578 2150 5590 2202
rect 5590 2150 5620 2202
rect 5644 2150 5654 2202
rect 5654 2150 5700 2202
rect 5404 2148 5460 2150
rect 5484 2148 5540 2150
rect 5564 2148 5620 2150
rect 5644 2148 5700 2150
rect 9852 2202 9908 2204
rect 9932 2202 9988 2204
rect 10012 2202 10068 2204
rect 10092 2202 10148 2204
rect 9852 2150 9898 2202
rect 9898 2150 9908 2202
rect 9932 2150 9962 2202
rect 9962 2150 9974 2202
rect 9974 2150 9988 2202
rect 10012 2150 10026 2202
rect 10026 2150 10038 2202
rect 10038 2150 10068 2202
rect 10092 2150 10102 2202
rect 10102 2150 10148 2202
rect 9852 2148 9908 2150
rect 9932 2148 9988 2150
rect 10012 2148 10068 2150
rect 10092 2148 10148 2150
rect 14300 2202 14356 2204
rect 14380 2202 14436 2204
rect 14460 2202 14516 2204
rect 14540 2202 14596 2204
rect 14300 2150 14346 2202
rect 14346 2150 14356 2202
rect 14380 2150 14410 2202
rect 14410 2150 14422 2202
rect 14422 2150 14436 2202
rect 14460 2150 14474 2202
rect 14474 2150 14486 2202
rect 14486 2150 14516 2202
rect 14540 2150 14550 2202
rect 14550 2150 14596 2202
rect 14300 2148 14356 2150
rect 14380 2148 14436 2150
rect 14460 2148 14516 2150
rect 14540 2148 14596 2150
<< metal3 >>
rect 5394 17440 5710 17441
rect 5394 17376 5400 17440
rect 5464 17376 5480 17440
rect 5544 17376 5560 17440
rect 5624 17376 5640 17440
rect 5704 17376 5710 17440
rect 5394 17375 5710 17376
rect 9842 17440 10158 17441
rect 9842 17376 9848 17440
rect 9912 17376 9928 17440
rect 9992 17376 10008 17440
rect 10072 17376 10088 17440
rect 10152 17376 10158 17440
rect 9842 17375 10158 17376
rect 14290 17440 14606 17441
rect 14290 17376 14296 17440
rect 14360 17376 14376 17440
rect 14440 17376 14456 17440
rect 14520 17376 14536 17440
rect 14600 17376 14606 17440
rect 14290 17375 14606 17376
rect 3170 16896 3486 16897
rect 3170 16832 3176 16896
rect 3240 16832 3256 16896
rect 3320 16832 3336 16896
rect 3400 16832 3416 16896
rect 3480 16832 3486 16896
rect 3170 16831 3486 16832
rect 7618 16896 7934 16897
rect 7618 16832 7624 16896
rect 7688 16832 7704 16896
rect 7768 16832 7784 16896
rect 7848 16832 7864 16896
rect 7928 16832 7934 16896
rect 7618 16831 7934 16832
rect 12066 16896 12382 16897
rect 12066 16832 12072 16896
rect 12136 16832 12152 16896
rect 12216 16832 12232 16896
rect 12296 16832 12312 16896
rect 12376 16832 12382 16896
rect 12066 16831 12382 16832
rect 16514 16896 16830 16897
rect 16514 16832 16520 16896
rect 16584 16832 16600 16896
rect 16664 16832 16680 16896
rect 16744 16832 16760 16896
rect 16824 16832 16830 16896
rect 16514 16831 16830 16832
rect 0 16418 800 16448
rect 1393 16418 1459 16421
rect 0 16416 1459 16418
rect 0 16360 1398 16416
rect 1454 16360 1459 16416
rect 0 16358 1459 16360
rect 0 16328 800 16358
rect 1393 16355 1459 16358
rect 5394 16352 5710 16353
rect 5394 16288 5400 16352
rect 5464 16288 5480 16352
rect 5544 16288 5560 16352
rect 5624 16288 5640 16352
rect 5704 16288 5710 16352
rect 5394 16287 5710 16288
rect 9842 16352 10158 16353
rect 9842 16288 9848 16352
rect 9912 16288 9928 16352
rect 9992 16288 10008 16352
rect 10072 16288 10088 16352
rect 10152 16288 10158 16352
rect 9842 16287 10158 16288
rect 14290 16352 14606 16353
rect 14290 16288 14296 16352
rect 14360 16288 14376 16352
rect 14440 16288 14456 16352
rect 14520 16288 14536 16352
rect 14600 16288 14606 16352
rect 14290 16287 14606 16288
rect 3170 15808 3486 15809
rect 3170 15744 3176 15808
rect 3240 15744 3256 15808
rect 3320 15744 3336 15808
rect 3400 15744 3416 15808
rect 3480 15744 3486 15808
rect 3170 15743 3486 15744
rect 7618 15808 7934 15809
rect 7618 15744 7624 15808
rect 7688 15744 7704 15808
rect 7768 15744 7784 15808
rect 7848 15744 7864 15808
rect 7928 15744 7934 15808
rect 7618 15743 7934 15744
rect 12066 15808 12382 15809
rect 12066 15744 12072 15808
rect 12136 15744 12152 15808
rect 12216 15744 12232 15808
rect 12296 15744 12312 15808
rect 12376 15744 12382 15808
rect 12066 15743 12382 15744
rect 16514 15808 16830 15809
rect 16514 15744 16520 15808
rect 16584 15744 16600 15808
rect 16664 15744 16680 15808
rect 16744 15744 16760 15808
rect 16824 15744 16830 15808
rect 16514 15743 16830 15744
rect 5394 15264 5710 15265
rect 5394 15200 5400 15264
rect 5464 15200 5480 15264
rect 5544 15200 5560 15264
rect 5624 15200 5640 15264
rect 5704 15200 5710 15264
rect 5394 15199 5710 15200
rect 9842 15264 10158 15265
rect 9842 15200 9848 15264
rect 9912 15200 9928 15264
rect 9992 15200 10008 15264
rect 10072 15200 10088 15264
rect 10152 15200 10158 15264
rect 9842 15199 10158 15200
rect 14290 15264 14606 15265
rect 14290 15200 14296 15264
rect 14360 15200 14376 15264
rect 14440 15200 14456 15264
rect 14520 15200 14536 15264
rect 14600 15200 14606 15264
rect 14290 15199 14606 15200
rect 3170 14720 3486 14721
rect 3170 14656 3176 14720
rect 3240 14656 3256 14720
rect 3320 14656 3336 14720
rect 3400 14656 3416 14720
rect 3480 14656 3486 14720
rect 3170 14655 3486 14656
rect 7618 14720 7934 14721
rect 7618 14656 7624 14720
rect 7688 14656 7704 14720
rect 7768 14656 7784 14720
rect 7848 14656 7864 14720
rect 7928 14656 7934 14720
rect 7618 14655 7934 14656
rect 12066 14720 12382 14721
rect 12066 14656 12072 14720
rect 12136 14656 12152 14720
rect 12216 14656 12232 14720
rect 12296 14656 12312 14720
rect 12376 14656 12382 14720
rect 12066 14655 12382 14656
rect 16514 14720 16830 14721
rect 16514 14656 16520 14720
rect 16584 14656 16600 14720
rect 16664 14656 16680 14720
rect 16744 14656 16760 14720
rect 16824 14656 16830 14720
rect 16514 14655 16830 14656
rect 5394 14176 5710 14177
rect 5394 14112 5400 14176
rect 5464 14112 5480 14176
rect 5544 14112 5560 14176
rect 5624 14112 5640 14176
rect 5704 14112 5710 14176
rect 5394 14111 5710 14112
rect 9842 14176 10158 14177
rect 9842 14112 9848 14176
rect 9912 14112 9928 14176
rect 9992 14112 10008 14176
rect 10072 14112 10088 14176
rect 10152 14112 10158 14176
rect 9842 14111 10158 14112
rect 14290 14176 14606 14177
rect 14290 14112 14296 14176
rect 14360 14112 14376 14176
rect 14440 14112 14456 14176
rect 14520 14112 14536 14176
rect 14600 14112 14606 14176
rect 14290 14111 14606 14112
rect 3170 13632 3486 13633
rect 3170 13568 3176 13632
rect 3240 13568 3256 13632
rect 3320 13568 3336 13632
rect 3400 13568 3416 13632
rect 3480 13568 3486 13632
rect 3170 13567 3486 13568
rect 7618 13632 7934 13633
rect 7618 13568 7624 13632
rect 7688 13568 7704 13632
rect 7768 13568 7784 13632
rect 7848 13568 7864 13632
rect 7928 13568 7934 13632
rect 7618 13567 7934 13568
rect 12066 13632 12382 13633
rect 12066 13568 12072 13632
rect 12136 13568 12152 13632
rect 12216 13568 12232 13632
rect 12296 13568 12312 13632
rect 12376 13568 12382 13632
rect 12066 13567 12382 13568
rect 16514 13632 16830 13633
rect 16514 13568 16520 13632
rect 16584 13568 16600 13632
rect 16664 13568 16680 13632
rect 16744 13568 16760 13632
rect 16824 13568 16830 13632
rect 16514 13567 16830 13568
rect 5394 13088 5710 13089
rect 5394 13024 5400 13088
rect 5464 13024 5480 13088
rect 5544 13024 5560 13088
rect 5624 13024 5640 13088
rect 5704 13024 5710 13088
rect 5394 13023 5710 13024
rect 9842 13088 10158 13089
rect 9842 13024 9848 13088
rect 9912 13024 9928 13088
rect 9992 13024 10008 13088
rect 10072 13024 10088 13088
rect 10152 13024 10158 13088
rect 9842 13023 10158 13024
rect 14290 13088 14606 13089
rect 14290 13024 14296 13088
rect 14360 13024 14376 13088
rect 14440 13024 14456 13088
rect 14520 13024 14536 13088
rect 14600 13024 14606 13088
rect 14290 13023 14606 13024
rect 3170 12544 3486 12545
rect 3170 12480 3176 12544
rect 3240 12480 3256 12544
rect 3320 12480 3336 12544
rect 3400 12480 3416 12544
rect 3480 12480 3486 12544
rect 3170 12479 3486 12480
rect 7618 12544 7934 12545
rect 7618 12480 7624 12544
rect 7688 12480 7704 12544
rect 7768 12480 7784 12544
rect 7848 12480 7864 12544
rect 7928 12480 7934 12544
rect 7618 12479 7934 12480
rect 12066 12544 12382 12545
rect 12066 12480 12072 12544
rect 12136 12480 12152 12544
rect 12216 12480 12232 12544
rect 12296 12480 12312 12544
rect 12376 12480 12382 12544
rect 12066 12479 12382 12480
rect 16514 12544 16830 12545
rect 16514 12480 16520 12544
rect 16584 12480 16600 12544
rect 16664 12480 16680 12544
rect 16744 12480 16760 12544
rect 16824 12480 16830 12544
rect 16514 12479 16830 12480
rect 5394 12000 5710 12001
rect 5394 11936 5400 12000
rect 5464 11936 5480 12000
rect 5544 11936 5560 12000
rect 5624 11936 5640 12000
rect 5704 11936 5710 12000
rect 5394 11935 5710 11936
rect 9842 12000 10158 12001
rect 9842 11936 9848 12000
rect 9912 11936 9928 12000
rect 9992 11936 10008 12000
rect 10072 11936 10088 12000
rect 10152 11936 10158 12000
rect 9842 11935 10158 11936
rect 14290 12000 14606 12001
rect 14290 11936 14296 12000
rect 14360 11936 14376 12000
rect 14440 11936 14456 12000
rect 14520 11936 14536 12000
rect 14600 11936 14606 12000
rect 14290 11935 14606 11936
rect 18137 11658 18203 11661
rect 19200 11658 20000 11688
rect 18137 11656 20000 11658
rect 18137 11600 18142 11656
rect 18198 11600 20000 11656
rect 18137 11598 20000 11600
rect 18137 11595 18203 11598
rect 19200 11568 20000 11598
rect 3170 11456 3486 11457
rect 3170 11392 3176 11456
rect 3240 11392 3256 11456
rect 3320 11392 3336 11456
rect 3400 11392 3416 11456
rect 3480 11392 3486 11456
rect 3170 11391 3486 11392
rect 7618 11456 7934 11457
rect 7618 11392 7624 11456
rect 7688 11392 7704 11456
rect 7768 11392 7784 11456
rect 7848 11392 7864 11456
rect 7928 11392 7934 11456
rect 7618 11391 7934 11392
rect 12066 11456 12382 11457
rect 12066 11392 12072 11456
rect 12136 11392 12152 11456
rect 12216 11392 12232 11456
rect 12296 11392 12312 11456
rect 12376 11392 12382 11456
rect 12066 11391 12382 11392
rect 16514 11456 16830 11457
rect 16514 11392 16520 11456
rect 16584 11392 16600 11456
rect 16664 11392 16680 11456
rect 16744 11392 16760 11456
rect 16824 11392 16830 11456
rect 16514 11391 16830 11392
rect 5394 10912 5710 10913
rect 5394 10848 5400 10912
rect 5464 10848 5480 10912
rect 5544 10848 5560 10912
rect 5624 10848 5640 10912
rect 5704 10848 5710 10912
rect 5394 10847 5710 10848
rect 9842 10912 10158 10913
rect 9842 10848 9848 10912
rect 9912 10848 9928 10912
rect 9992 10848 10008 10912
rect 10072 10848 10088 10912
rect 10152 10848 10158 10912
rect 9842 10847 10158 10848
rect 14290 10912 14606 10913
rect 14290 10848 14296 10912
rect 14360 10848 14376 10912
rect 14440 10848 14456 10912
rect 14520 10848 14536 10912
rect 14600 10848 14606 10912
rect 14290 10847 14606 10848
rect 3170 10368 3486 10369
rect 3170 10304 3176 10368
rect 3240 10304 3256 10368
rect 3320 10304 3336 10368
rect 3400 10304 3416 10368
rect 3480 10304 3486 10368
rect 3170 10303 3486 10304
rect 7618 10368 7934 10369
rect 7618 10304 7624 10368
rect 7688 10304 7704 10368
rect 7768 10304 7784 10368
rect 7848 10304 7864 10368
rect 7928 10304 7934 10368
rect 7618 10303 7934 10304
rect 12066 10368 12382 10369
rect 12066 10304 12072 10368
rect 12136 10304 12152 10368
rect 12216 10304 12232 10368
rect 12296 10304 12312 10368
rect 12376 10304 12382 10368
rect 12066 10303 12382 10304
rect 16514 10368 16830 10369
rect 16514 10304 16520 10368
rect 16584 10304 16600 10368
rect 16664 10304 16680 10368
rect 16744 10304 16760 10368
rect 16824 10304 16830 10368
rect 16514 10303 16830 10304
rect 5394 9824 5710 9825
rect 5394 9760 5400 9824
rect 5464 9760 5480 9824
rect 5544 9760 5560 9824
rect 5624 9760 5640 9824
rect 5704 9760 5710 9824
rect 5394 9759 5710 9760
rect 9842 9824 10158 9825
rect 9842 9760 9848 9824
rect 9912 9760 9928 9824
rect 9992 9760 10008 9824
rect 10072 9760 10088 9824
rect 10152 9760 10158 9824
rect 9842 9759 10158 9760
rect 14290 9824 14606 9825
rect 14290 9760 14296 9824
rect 14360 9760 14376 9824
rect 14440 9760 14456 9824
rect 14520 9760 14536 9824
rect 14600 9760 14606 9824
rect 14290 9759 14606 9760
rect 3170 9280 3486 9281
rect 3170 9216 3176 9280
rect 3240 9216 3256 9280
rect 3320 9216 3336 9280
rect 3400 9216 3416 9280
rect 3480 9216 3486 9280
rect 3170 9215 3486 9216
rect 7618 9280 7934 9281
rect 7618 9216 7624 9280
rect 7688 9216 7704 9280
rect 7768 9216 7784 9280
rect 7848 9216 7864 9280
rect 7928 9216 7934 9280
rect 7618 9215 7934 9216
rect 12066 9280 12382 9281
rect 12066 9216 12072 9280
rect 12136 9216 12152 9280
rect 12216 9216 12232 9280
rect 12296 9216 12312 9280
rect 12376 9216 12382 9280
rect 12066 9215 12382 9216
rect 16514 9280 16830 9281
rect 16514 9216 16520 9280
rect 16584 9216 16600 9280
rect 16664 9216 16680 9280
rect 16744 9216 16760 9280
rect 16824 9216 16830 9280
rect 16514 9215 16830 9216
rect 5394 8736 5710 8737
rect 5394 8672 5400 8736
rect 5464 8672 5480 8736
rect 5544 8672 5560 8736
rect 5624 8672 5640 8736
rect 5704 8672 5710 8736
rect 5394 8671 5710 8672
rect 9842 8736 10158 8737
rect 9842 8672 9848 8736
rect 9912 8672 9928 8736
rect 9992 8672 10008 8736
rect 10072 8672 10088 8736
rect 10152 8672 10158 8736
rect 9842 8671 10158 8672
rect 14290 8736 14606 8737
rect 14290 8672 14296 8736
rect 14360 8672 14376 8736
rect 14440 8672 14456 8736
rect 14520 8672 14536 8736
rect 14600 8672 14606 8736
rect 14290 8671 14606 8672
rect 3170 8192 3486 8193
rect 3170 8128 3176 8192
rect 3240 8128 3256 8192
rect 3320 8128 3336 8192
rect 3400 8128 3416 8192
rect 3480 8128 3486 8192
rect 3170 8127 3486 8128
rect 7618 8192 7934 8193
rect 7618 8128 7624 8192
rect 7688 8128 7704 8192
rect 7768 8128 7784 8192
rect 7848 8128 7864 8192
rect 7928 8128 7934 8192
rect 7618 8127 7934 8128
rect 12066 8192 12382 8193
rect 12066 8128 12072 8192
rect 12136 8128 12152 8192
rect 12216 8128 12232 8192
rect 12296 8128 12312 8192
rect 12376 8128 12382 8192
rect 12066 8127 12382 8128
rect 16514 8192 16830 8193
rect 16514 8128 16520 8192
rect 16584 8128 16600 8192
rect 16664 8128 16680 8192
rect 16744 8128 16760 8192
rect 16824 8128 16830 8192
rect 16514 8127 16830 8128
rect 5394 7648 5710 7649
rect 5394 7584 5400 7648
rect 5464 7584 5480 7648
rect 5544 7584 5560 7648
rect 5624 7584 5640 7648
rect 5704 7584 5710 7648
rect 5394 7583 5710 7584
rect 9842 7648 10158 7649
rect 9842 7584 9848 7648
rect 9912 7584 9928 7648
rect 9992 7584 10008 7648
rect 10072 7584 10088 7648
rect 10152 7584 10158 7648
rect 9842 7583 10158 7584
rect 14290 7648 14606 7649
rect 14290 7584 14296 7648
rect 14360 7584 14376 7648
rect 14440 7584 14456 7648
rect 14520 7584 14536 7648
rect 14600 7584 14606 7648
rect 14290 7583 14606 7584
rect 3170 7104 3486 7105
rect 3170 7040 3176 7104
rect 3240 7040 3256 7104
rect 3320 7040 3336 7104
rect 3400 7040 3416 7104
rect 3480 7040 3486 7104
rect 3170 7039 3486 7040
rect 7618 7104 7934 7105
rect 7618 7040 7624 7104
rect 7688 7040 7704 7104
rect 7768 7040 7784 7104
rect 7848 7040 7864 7104
rect 7928 7040 7934 7104
rect 7618 7039 7934 7040
rect 12066 7104 12382 7105
rect 12066 7040 12072 7104
rect 12136 7040 12152 7104
rect 12216 7040 12232 7104
rect 12296 7040 12312 7104
rect 12376 7040 12382 7104
rect 12066 7039 12382 7040
rect 16514 7104 16830 7105
rect 16514 7040 16520 7104
rect 16584 7040 16600 7104
rect 16664 7040 16680 7104
rect 16744 7040 16760 7104
rect 16824 7040 16830 7104
rect 16514 7039 16830 7040
rect 5394 6560 5710 6561
rect 5394 6496 5400 6560
rect 5464 6496 5480 6560
rect 5544 6496 5560 6560
rect 5624 6496 5640 6560
rect 5704 6496 5710 6560
rect 5394 6495 5710 6496
rect 9842 6560 10158 6561
rect 9842 6496 9848 6560
rect 9912 6496 9928 6560
rect 9992 6496 10008 6560
rect 10072 6496 10088 6560
rect 10152 6496 10158 6560
rect 9842 6495 10158 6496
rect 14290 6560 14606 6561
rect 14290 6496 14296 6560
rect 14360 6496 14376 6560
rect 14440 6496 14456 6560
rect 14520 6496 14536 6560
rect 14600 6496 14606 6560
rect 14290 6495 14606 6496
rect 3170 6016 3486 6017
rect 3170 5952 3176 6016
rect 3240 5952 3256 6016
rect 3320 5952 3336 6016
rect 3400 5952 3416 6016
rect 3480 5952 3486 6016
rect 3170 5951 3486 5952
rect 7618 6016 7934 6017
rect 7618 5952 7624 6016
rect 7688 5952 7704 6016
rect 7768 5952 7784 6016
rect 7848 5952 7864 6016
rect 7928 5952 7934 6016
rect 7618 5951 7934 5952
rect 12066 6016 12382 6017
rect 12066 5952 12072 6016
rect 12136 5952 12152 6016
rect 12216 5952 12232 6016
rect 12296 5952 12312 6016
rect 12376 5952 12382 6016
rect 12066 5951 12382 5952
rect 16514 6016 16830 6017
rect 16514 5952 16520 6016
rect 16584 5952 16600 6016
rect 16664 5952 16680 6016
rect 16744 5952 16760 6016
rect 16824 5952 16830 6016
rect 16514 5951 16830 5952
rect 5394 5472 5710 5473
rect 5394 5408 5400 5472
rect 5464 5408 5480 5472
rect 5544 5408 5560 5472
rect 5624 5408 5640 5472
rect 5704 5408 5710 5472
rect 5394 5407 5710 5408
rect 9842 5472 10158 5473
rect 9842 5408 9848 5472
rect 9912 5408 9928 5472
rect 9992 5408 10008 5472
rect 10072 5408 10088 5472
rect 10152 5408 10158 5472
rect 9842 5407 10158 5408
rect 14290 5472 14606 5473
rect 14290 5408 14296 5472
rect 14360 5408 14376 5472
rect 14440 5408 14456 5472
rect 14520 5408 14536 5472
rect 14600 5408 14606 5472
rect 14290 5407 14606 5408
rect 3170 4928 3486 4929
rect 3170 4864 3176 4928
rect 3240 4864 3256 4928
rect 3320 4864 3336 4928
rect 3400 4864 3416 4928
rect 3480 4864 3486 4928
rect 3170 4863 3486 4864
rect 7618 4928 7934 4929
rect 7618 4864 7624 4928
rect 7688 4864 7704 4928
rect 7768 4864 7784 4928
rect 7848 4864 7864 4928
rect 7928 4864 7934 4928
rect 7618 4863 7934 4864
rect 12066 4928 12382 4929
rect 12066 4864 12072 4928
rect 12136 4864 12152 4928
rect 12216 4864 12232 4928
rect 12296 4864 12312 4928
rect 12376 4864 12382 4928
rect 12066 4863 12382 4864
rect 16514 4928 16830 4929
rect 16514 4864 16520 4928
rect 16584 4864 16600 4928
rect 16664 4864 16680 4928
rect 16744 4864 16760 4928
rect 16824 4864 16830 4928
rect 16514 4863 16830 4864
rect 5394 4384 5710 4385
rect 5394 4320 5400 4384
rect 5464 4320 5480 4384
rect 5544 4320 5560 4384
rect 5624 4320 5640 4384
rect 5704 4320 5710 4384
rect 5394 4319 5710 4320
rect 9842 4384 10158 4385
rect 9842 4320 9848 4384
rect 9912 4320 9928 4384
rect 9992 4320 10008 4384
rect 10072 4320 10088 4384
rect 10152 4320 10158 4384
rect 9842 4319 10158 4320
rect 14290 4384 14606 4385
rect 14290 4320 14296 4384
rect 14360 4320 14376 4384
rect 14440 4320 14456 4384
rect 14520 4320 14536 4384
rect 14600 4320 14606 4384
rect 14290 4319 14606 4320
rect 3170 3840 3486 3841
rect 3170 3776 3176 3840
rect 3240 3776 3256 3840
rect 3320 3776 3336 3840
rect 3400 3776 3416 3840
rect 3480 3776 3486 3840
rect 3170 3775 3486 3776
rect 7618 3840 7934 3841
rect 7618 3776 7624 3840
rect 7688 3776 7704 3840
rect 7768 3776 7784 3840
rect 7848 3776 7864 3840
rect 7928 3776 7934 3840
rect 7618 3775 7934 3776
rect 12066 3840 12382 3841
rect 12066 3776 12072 3840
rect 12136 3776 12152 3840
rect 12216 3776 12232 3840
rect 12296 3776 12312 3840
rect 12376 3776 12382 3840
rect 12066 3775 12382 3776
rect 16514 3840 16830 3841
rect 16514 3776 16520 3840
rect 16584 3776 16600 3840
rect 16664 3776 16680 3840
rect 16744 3776 16760 3840
rect 16824 3776 16830 3840
rect 16514 3775 16830 3776
rect 5394 3296 5710 3297
rect 5394 3232 5400 3296
rect 5464 3232 5480 3296
rect 5544 3232 5560 3296
rect 5624 3232 5640 3296
rect 5704 3232 5710 3296
rect 5394 3231 5710 3232
rect 9842 3296 10158 3297
rect 9842 3232 9848 3296
rect 9912 3232 9928 3296
rect 9992 3232 10008 3296
rect 10072 3232 10088 3296
rect 10152 3232 10158 3296
rect 9842 3231 10158 3232
rect 14290 3296 14606 3297
rect 14290 3232 14296 3296
rect 14360 3232 14376 3296
rect 14440 3232 14456 3296
rect 14520 3232 14536 3296
rect 14600 3232 14606 3296
rect 14290 3231 14606 3232
rect 3170 2752 3486 2753
rect 3170 2688 3176 2752
rect 3240 2688 3256 2752
rect 3320 2688 3336 2752
rect 3400 2688 3416 2752
rect 3480 2688 3486 2752
rect 3170 2687 3486 2688
rect 7618 2752 7934 2753
rect 7618 2688 7624 2752
rect 7688 2688 7704 2752
rect 7768 2688 7784 2752
rect 7848 2688 7864 2752
rect 7928 2688 7934 2752
rect 7618 2687 7934 2688
rect 12066 2752 12382 2753
rect 12066 2688 12072 2752
rect 12136 2688 12152 2752
rect 12216 2688 12232 2752
rect 12296 2688 12312 2752
rect 12376 2688 12382 2752
rect 12066 2687 12382 2688
rect 16514 2752 16830 2753
rect 16514 2688 16520 2752
rect 16584 2688 16600 2752
rect 16664 2688 16680 2752
rect 16744 2688 16760 2752
rect 16824 2688 16830 2752
rect 16514 2687 16830 2688
rect 5394 2208 5710 2209
rect 5394 2144 5400 2208
rect 5464 2144 5480 2208
rect 5544 2144 5560 2208
rect 5624 2144 5640 2208
rect 5704 2144 5710 2208
rect 5394 2143 5710 2144
rect 9842 2208 10158 2209
rect 9842 2144 9848 2208
rect 9912 2144 9928 2208
rect 9992 2144 10008 2208
rect 10072 2144 10088 2208
rect 10152 2144 10158 2208
rect 9842 2143 10158 2144
rect 14290 2208 14606 2209
rect 14290 2144 14296 2208
rect 14360 2144 14376 2208
rect 14440 2144 14456 2208
rect 14520 2144 14536 2208
rect 14600 2144 14606 2208
rect 14290 2143 14606 2144
<< via3 >>
rect 5400 17436 5464 17440
rect 5400 17380 5404 17436
rect 5404 17380 5460 17436
rect 5460 17380 5464 17436
rect 5400 17376 5464 17380
rect 5480 17436 5544 17440
rect 5480 17380 5484 17436
rect 5484 17380 5540 17436
rect 5540 17380 5544 17436
rect 5480 17376 5544 17380
rect 5560 17436 5624 17440
rect 5560 17380 5564 17436
rect 5564 17380 5620 17436
rect 5620 17380 5624 17436
rect 5560 17376 5624 17380
rect 5640 17436 5704 17440
rect 5640 17380 5644 17436
rect 5644 17380 5700 17436
rect 5700 17380 5704 17436
rect 5640 17376 5704 17380
rect 9848 17436 9912 17440
rect 9848 17380 9852 17436
rect 9852 17380 9908 17436
rect 9908 17380 9912 17436
rect 9848 17376 9912 17380
rect 9928 17436 9992 17440
rect 9928 17380 9932 17436
rect 9932 17380 9988 17436
rect 9988 17380 9992 17436
rect 9928 17376 9992 17380
rect 10008 17436 10072 17440
rect 10008 17380 10012 17436
rect 10012 17380 10068 17436
rect 10068 17380 10072 17436
rect 10008 17376 10072 17380
rect 10088 17436 10152 17440
rect 10088 17380 10092 17436
rect 10092 17380 10148 17436
rect 10148 17380 10152 17436
rect 10088 17376 10152 17380
rect 14296 17436 14360 17440
rect 14296 17380 14300 17436
rect 14300 17380 14356 17436
rect 14356 17380 14360 17436
rect 14296 17376 14360 17380
rect 14376 17436 14440 17440
rect 14376 17380 14380 17436
rect 14380 17380 14436 17436
rect 14436 17380 14440 17436
rect 14376 17376 14440 17380
rect 14456 17436 14520 17440
rect 14456 17380 14460 17436
rect 14460 17380 14516 17436
rect 14516 17380 14520 17436
rect 14456 17376 14520 17380
rect 14536 17436 14600 17440
rect 14536 17380 14540 17436
rect 14540 17380 14596 17436
rect 14596 17380 14600 17436
rect 14536 17376 14600 17380
rect 3176 16892 3240 16896
rect 3176 16836 3180 16892
rect 3180 16836 3236 16892
rect 3236 16836 3240 16892
rect 3176 16832 3240 16836
rect 3256 16892 3320 16896
rect 3256 16836 3260 16892
rect 3260 16836 3316 16892
rect 3316 16836 3320 16892
rect 3256 16832 3320 16836
rect 3336 16892 3400 16896
rect 3336 16836 3340 16892
rect 3340 16836 3396 16892
rect 3396 16836 3400 16892
rect 3336 16832 3400 16836
rect 3416 16892 3480 16896
rect 3416 16836 3420 16892
rect 3420 16836 3476 16892
rect 3476 16836 3480 16892
rect 3416 16832 3480 16836
rect 7624 16892 7688 16896
rect 7624 16836 7628 16892
rect 7628 16836 7684 16892
rect 7684 16836 7688 16892
rect 7624 16832 7688 16836
rect 7704 16892 7768 16896
rect 7704 16836 7708 16892
rect 7708 16836 7764 16892
rect 7764 16836 7768 16892
rect 7704 16832 7768 16836
rect 7784 16892 7848 16896
rect 7784 16836 7788 16892
rect 7788 16836 7844 16892
rect 7844 16836 7848 16892
rect 7784 16832 7848 16836
rect 7864 16892 7928 16896
rect 7864 16836 7868 16892
rect 7868 16836 7924 16892
rect 7924 16836 7928 16892
rect 7864 16832 7928 16836
rect 12072 16892 12136 16896
rect 12072 16836 12076 16892
rect 12076 16836 12132 16892
rect 12132 16836 12136 16892
rect 12072 16832 12136 16836
rect 12152 16892 12216 16896
rect 12152 16836 12156 16892
rect 12156 16836 12212 16892
rect 12212 16836 12216 16892
rect 12152 16832 12216 16836
rect 12232 16892 12296 16896
rect 12232 16836 12236 16892
rect 12236 16836 12292 16892
rect 12292 16836 12296 16892
rect 12232 16832 12296 16836
rect 12312 16892 12376 16896
rect 12312 16836 12316 16892
rect 12316 16836 12372 16892
rect 12372 16836 12376 16892
rect 12312 16832 12376 16836
rect 16520 16892 16584 16896
rect 16520 16836 16524 16892
rect 16524 16836 16580 16892
rect 16580 16836 16584 16892
rect 16520 16832 16584 16836
rect 16600 16892 16664 16896
rect 16600 16836 16604 16892
rect 16604 16836 16660 16892
rect 16660 16836 16664 16892
rect 16600 16832 16664 16836
rect 16680 16892 16744 16896
rect 16680 16836 16684 16892
rect 16684 16836 16740 16892
rect 16740 16836 16744 16892
rect 16680 16832 16744 16836
rect 16760 16892 16824 16896
rect 16760 16836 16764 16892
rect 16764 16836 16820 16892
rect 16820 16836 16824 16892
rect 16760 16832 16824 16836
rect 5400 16348 5464 16352
rect 5400 16292 5404 16348
rect 5404 16292 5460 16348
rect 5460 16292 5464 16348
rect 5400 16288 5464 16292
rect 5480 16348 5544 16352
rect 5480 16292 5484 16348
rect 5484 16292 5540 16348
rect 5540 16292 5544 16348
rect 5480 16288 5544 16292
rect 5560 16348 5624 16352
rect 5560 16292 5564 16348
rect 5564 16292 5620 16348
rect 5620 16292 5624 16348
rect 5560 16288 5624 16292
rect 5640 16348 5704 16352
rect 5640 16292 5644 16348
rect 5644 16292 5700 16348
rect 5700 16292 5704 16348
rect 5640 16288 5704 16292
rect 9848 16348 9912 16352
rect 9848 16292 9852 16348
rect 9852 16292 9908 16348
rect 9908 16292 9912 16348
rect 9848 16288 9912 16292
rect 9928 16348 9992 16352
rect 9928 16292 9932 16348
rect 9932 16292 9988 16348
rect 9988 16292 9992 16348
rect 9928 16288 9992 16292
rect 10008 16348 10072 16352
rect 10008 16292 10012 16348
rect 10012 16292 10068 16348
rect 10068 16292 10072 16348
rect 10008 16288 10072 16292
rect 10088 16348 10152 16352
rect 10088 16292 10092 16348
rect 10092 16292 10148 16348
rect 10148 16292 10152 16348
rect 10088 16288 10152 16292
rect 14296 16348 14360 16352
rect 14296 16292 14300 16348
rect 14300 16292 14356 16348
rect 14356 16292 14360 16348
rect 14296 16288 14360 16292
rect 14376 16348 14440 16352
rect 14376 16292 14380 16348
rect 14380 16292 14436 16348
rect 14436 16292 14440 16348
rect 14376 16288 14440 16292
rect 14456 16348 14520 16352
rect 14456 16292 14460 16348
rect 14460 16292 14516 16348
rect 14516 16292 14520 16348
rect 14456 16288 14520 16292
rect 14536 16348 14600 16352
rect 14536 16292 14540 16348
rect 14540 16292 14596 16348
rect 14596 16292 14600 16348
rect 14536 16288 14600 16292
rect 3176 15804 3240 15808
rect 3176 15748 3180 15804
rect 3180 15748 3236 15804
rect 3236 15748 3240 15804
rect 3176 15744 3240 15748
rect 3256 15804 3320 15808
rect 3256 15748 3260 15804
rect 3260 15748 3316 15804
rect 3316 15748 3320 15804
rect 3256 15744 3320 15748
rect 3336 15804 3400 15808
rect 3336 15748 3340 15804
rect 3340 15748 3396 15804
rect 3396 15748 3400 15804
rect 3336 15744 3400 15748
rect 3416 15804 3480 15808
rect 3416 15748 3420 15804
rect 3420 15748 3476 15804
rect 3476 15748 3480 15804
rect 3416 15744 3480 15748
rect 7624 15804 7688 15808
rect 7624 15748 7628 15804
rect 7628 15748 7684 15804
rect 7684 15748 7688 15804
rect 7624 15744 7688 15748
rect 7704 15804 7768 15808
rect 7704 15748 7708 15804
rect 7708 15748 7764 15804
rect 7764 15748 7768 15804
rect 7704 15744 7768 15748
rect 7784 15804 7848 15808
rect 7784 15748 7788 15804
rect 7788 15748 7844 15804
rect 7844 15748 7848 15804
rect 7784 15744 7848 15748
rect 7864 15804 7928 15808
rect 7864 15748 7868 15804
rect 7868 15748 7924 15804
rect 7924 15748 7928 15804
rect 7864 15744 7928 15748
rect 12072 15804 12136 15808
rect 12072 15748 12076 15804
rect 12076 15748 12132 15804
rect 12132 15748 12136 15804
rect 12072 15744 12136 15748
rect 12152 15804 12216 15808
rect 12152 15748 12156 15804
rect 12156 15748 12212 15804
rect 12212 15748 12216 15804
rect 12152 15744 12216 15748
rect 12232 15804 12296 15808
rect 12232 15748 12236 15804
rect 12236 15748 12292 15804
rect 12292 15748 12296 15804
rect 12232 15744 12296 15748
rect 12312 15804 12376 15808
rect 12312 15748 12316 15804
rect 12316 15748 12372 15804
rect 12372 15748 12376 15804
rect 12312 15744 12376 15748
rect 16520 15804 16584 15808
rect 16520 15748 16524 15804
rect 16524 15748 16580 15804
rect 16580 15748 16584 15804
rect 16520 15744 16584 15748
rect 16600 15804 16664 15808
rect 16600 15748 16604 15804
rect 16604 15748 16660 15804
rect 16660 15748 16664 15804
rect 16600 15744 16664 15748
rect 16680 15804 16744 15808
rect 16680 15748 16684 15804
rect 16684 15748 16740 15804
rect 16740 15748 16744 15804
rect 16680 15744 16744 15748
rect 16760 15804 16824 15808
rect 16760 15748 16764 15804
rect 16764 15748 16820 15804
rect 16820 15748 16824 15804
rect 16760 15744 16824 15748
rect 5400 15260 5464 15264
rect 5400 15204 5404 15260
rect 5404 15204 5460 15260
rect 5460 15204 5464 15260
rect 5400 15200 5464 15204
rect 5480 15260 5544 15264
rect 5480 15204 5484 15260
rect 5484 15204 5540 15260
rect 5540 15204 5544 15260
rect 5480 15200 5544 15204
rect 5560 15260 5624 15264
rect 5560 15204 5564 15260
rect 5564 15204 5620 15260
rect 5620 15204 5624 15260
rect 5560 15200 5624 15204
rect 5640 15260 5704 15264
rect 5640 15204 5644 15260
rect 5644 15204 5700 15260
rect 5700 15204 5704 15260
rect 5640 15200 5704 15204
rect 9848 15260 9912 15264
rect 9848 15204 9852 15260
rect 9852 15204 9908 15260
rect 9908 15204 9912 15260
rect 9848 15200 9912 15204
rect 9928 15260 9992 15264
rect 9928 15204 9932 15260
rect 9932 15204 9988 15260
rect 9988 15204 9992 15260
rect 9928 15200 9992 15204
rect 10008 15260 10072 15264
rect 10008 15204 10012 15260
rect 10012 15204 10068 15260
rect 10068 15204 10072 15260
rect 10008 15200 10072 15204
rect 10088 15260 10152 15264
rect 10088 15204 10092 15260
rect 10092 15204 10148 15260
rect 10148 15204 10152 15260
rect 10088 15200 10152 15204
rect 14296 15260 14360 15264
rect 14296 15204 14300 15260
rect 14300 15204 14356 15260
rect 14356 15204 14360 15260
rect 14296 15200 14360 15204
rect 14376 15260 14440 15264
rect 14376 15204 14380 15260
rect 14380 15204 14436 15260
rect 14436 15204 14440 15260
rect 14376 15200 14440 15204
rect 14456 15260 14520 15264
rect 14456 15204 14460 15260
rect 14460 15204 14516 15260
rect 14516 15204 14520 15260
rect 14456 15200 14520 15204
rect 14536 15260 14600 15264
rect 14536 15204 14540 15260
rect 14540 15204 14596 15260
rect 14596 15204 14600 15260
rect 14536 15200 14600 15204
rect 3176 14716 3240 14720
rect 3176 14660 3180 14716
rect 3180 14660 3236 14716
rect 3236 14660 3240 14716
rect 3176 14656 3240 14660
rect 3256 14716 3320 14720
rect 3256 14660 3260 14716
rect 3260 14660 3316 14716
rect 3316 14660 3320 14716
rect 3256 14656 3320 14660
rect 3336 14716 3400 14720
rect 3336 14660 3340 14716
rect 3340 14660 3396 14716
rect 3396 14660 3400 14716
rect 3336 14656 3400 14660
rect 3416 14716 3480 14720
rect 3416 14660 3420 14716
rect 3420 14660 3476 14716
rect 3476 14660 3480 14716
rect 3416 14656 3480 14660
rect 7624 14716 7688 14720
rect 7624 14660 7628 14716
rect 7628 14660 7684 14716
rect 7684 14660 7688 14716
rect 7624 14656 7688 14660
rect 7704 14716 7768 14720
rect 7704 14660 7708 14716
rect 7708 14660 7764 14716
rect 7764 14660 7768 14716
rect 7704 14656 7768 14660
rect 7784 14716 7848 14720
rect 7784 14660 7788 14716
rect 7788 14660 7844 14716
rect 7844 14660 7848 14716
rect 7784 14656 7848 14660
rect 7864 14716 7928 14720
rect 7864 14660 7868 14716
rect 7868 14660 7924 14716
rect 7924 14660 7928 14716
rect 7864 14656 7928 14660
rect 12072 14716 12136 14720
rect 12072 14660 12076 14716
rect 12076 14660 12132 14716
rect 12132 14660 12136 14716
rect 12072 14656 12136 14660
rect 12152 14716 12216 14720
rect 12152 14660 12156 14716
rect 12156 14660 12212 14716
rect 12212 14660 12216 14716
rect 12152 14656 12216 14660
rect 12232 14716 12296 14720
rect 12232 14660 12236 14716
rect 12236 14660 12292 14716
rect 12292 14660 12296 14716
rect 12232 14656 12296 14660
rect 12312 14716 12376 14720
rect 12312 14660 12316 14716
rect 12316 14660 12372 14716
rect 12372 14660 12376 14716
rect 12312 14656 12376 14660
rect 16520 14716 16584 14720
rect 16520 14660 16524 14716
rect 16524 14660 16580 14716
rect 16580 14660 16584 14716
rect 16520 14656 16584 14660
rect 16600 14716 16664 14720
rect 16600 14660 16604 14716
rect 16604 14660 16660 14716
rect 16660 14660 16664 14716
rect 16600 14656 16664 14660
rect 16680 14716 16744 14720
rect 16680 14660 16684 14716
rect 16684 14660 16740 14716
rect 16740 14660 16744 14716
rect 16680 14656 16744 14660
rect 16760 14716 16824 14720
rect 16760 14660 16764 14716
rect 16764 14660 16820 14716
rect 16820 14660 16824 14716
rect 16760 14656 16824 14660
rect 5400 14172 5464 14176
rect 5400 14116 5404 14172
rect 5404 14116 5460 14172
rect 5460 14116 5464 14172
rect 5400 14112 5464 14116
rect 5480 14172 5544 14176
rect 5480 14116 5484 14172
rect 5484 14116 5540 14172
rect 5540 14116 5544 14172
rect 5480 14112 5544 14116
rect 5560 14172 5624 14176
rect 5560 14116 5564 14172
rect 5564 14116 5620 14172
rect 5620 14116 5624 14172
rect 5560 14112 5624 14116
rect 5640 14172 5704 14176
rect 5640 14116 5644 14172
rect 5644 14116 5700 14172
rect 5700 14116 5704 14172
rect 5640 14112 5704 14116
rect 9848 14172 9912 14176
rect 9848 14116 9852 14172
rect 9852 14116 9908 14172
rect 9908 14116 9912 14172
rect 9848 14112 9912 14116
rect 9928 14172 9992 14176
rect 9928 14116 9932 14172
rect 9932 14116 9988 14172
rect 9988 14116 9992 14172
rect 9928 14112 9992 14116
rect 10008 14172 10072 14176
rect 10008 14116 10012 14172
rect 10012 14116 10068 14172
rect 10068 14116 10072 14172
rect 10008 14112 10072 14116
rect 10088 14172 10152 14176
rect 10088 14116 10092 14172
rect 10092 14116 10148 14172
rect 10148 14116 10152 14172
rect 10088 14112 10152 14116
rect 14296 14172 14360 14176
rect 14296 14116 14300 14172
rect 14300 14116 14356 14172
rect 14356 14116 14360 14172
rect 14296 14112 14360 14116
rect 14376 14172 14440 14176
rect 14376 14116 14380 14172
rect 14380 14116 14436 14172
rect 14436 14116 14440 14172
rect 14376 14112 14440 14116
rect 14456 14172 14520 14176
rect 14456 14116 14460 14172
rect 14460 14116 14516 14172
rect 14516 14116 14520 14172
rect 14456 14112 14520 14116
rect 14536 14172 14600 14176
rect 14536 14116 14540 14172
rect 14540 14116 14596 14172
rect 14596 14116 14600 14172
rect 14536 14112 14600 14116
rect 3176 13628 3240 13632
rect 3176 13572 3180 13628
rect 3180 13572 3236 13628
rect 3236 13572 3240 13628
rect 3176 13568 3240 13572
rect 3256 13628 3320 13632
rect 3256 13572 3260 13628
rect 3260 13572 3316 13628
rect 3316 13572 3320 13628
rect 3256 13568 3320 13572
rect 3336 13628 3400 13632
rect 3336 13572 3340 13628
rect 3340 13572 3396 13628
rect 3396 13572 3400 13628
rect 3336 13568 3400 13572
rect 3416 13628 3480 13632
rect 3416 13572 3420 13628
rect 3420 13572 3476 13628
rect 3476 13572 3480 13628
rect 3416 13568 3480 13572
rect 7624 13628 7688 13632
rect 7624 13572 7628 13628
rect 7628 13572 7684 13628
rect 7684 13572 7688 13628
rect 7624 13568 7688 13572
rect 7704 13628 7768 13632
rect 7704 13572 7708 13628
rect 7708 13572 7764 13628
rect 7764 13572 7768 13628
rect 7704 13568 7768 13572
rect 7784 13628 7848 13632
rect 7784 13572 7788 13628
rect 7788 13572 7844 13628
rect 7844 13572 7848 13628
rect 7784 13568 7848 13572
rect 7864 13628 7928 13632
rect 7864 13572 7868 13628
rect 7868 13572 7924 13628
rect 7924 13572 7928 13628
rect 7864 13568 7928 13572
rect 12072 13628 12136 13632
rect 12072 13572 12076 13628
rect 12076 13572 12132 13628
rect 12132 13572 12136 13628
rect 12072 13568 12136 13572
rect 12152 13628 12216 13632
rect 12152 13572 12156 13628
rect 12156 13572 12212 13628
rect 12212 13572 12216 13628
rect 12152 13568 12216 13572
rect 12232 13628 12296 13632
rect 12232 13572 12236 13628
rect 12236 13572 12292 13628
rect 12292 13572 12296 13628
rect 12232 13568 12296 13572
rect 12312 13628 12376 13632
rect 12312 13572 12316 13628
rect 12316 13572 12372 13628
rect 12372 13572 12376 13628
rect 12312 13568 12376 13572
rect 16520 13628 16584 13632
rect 16520 13572 16524 13628
rect 16524 13572 16580 13628
rect 16580 13572 16584 13628
rect 16520 13568 16584 13572
rect 16600 13628 16664 13632
rect 16600 13572 16604 13628
rect 16604 13572 16660 13628
rect 16660 13572 16664 13628
rect 16600 13568 16664 13572
rect 16680 13628 16744 13632
rect 16680 13572 16684 13628
rect 16684 13572 16740 13628
rect 16740 13572 16744 13628
rect 16680 13568 16744 13572
rect 16760 13628 16824 13632
rect 16760 13572 16764 13628
rect 16764 13572 16820 13628
rect 16820 13572 16824 13628
rect 16760 13568 16824 13572
rect 5400 13084 5464 13088
rect 5400 13028 5404 13084
rect 5404 13028 5460 13084
rect 5460 13028 5464 13084
rect 5400 13024 5464 13028
rect 5480 13084 5544 13088
rect 5480 13028 5484 13084
rect 5484 13028 5540 13084
rect 5540 13028 5544 13084
rect 5480 13024 5544 13028
rect 5560 13084 5624 13088
rect 5560 13028 5564 13084
rect 5564 13028 5620 13084
rect 5620 13028 5624 13084
rect 5560 13024 5624 13028
rect 5640 13084 5704 13088
rect 5640 13028 5644 13084
rect 5644 13028 5700 13084
rect 5700 13028 5704 13084
rect 5640 13024 5704 13028
rect 9848 13084 9912 13088
rect 9848 13028 9852 13084
rect 9852 13028 9908 13084
rect 9908 13028 9912 13084
rect 9848 13024 9912 13028
rect 9928 13084 9992 13088
rect 9928 13028 9932 13084
rect 9932 13028 9988 13084
rect 9988 13028 9992 13084
rect 9928 13024 9992 13028
rect 10008 13084 10072 13088
rect 10008 13028 10012 13084
rect 10012 13028 10068 13084
rect 10068 13028 10072 13084
rect 10008 13024 10072 13028
rect 10088 13084 10152 13088
rect 10088 13028 10092 13084
rect 10092 13028 10148 13084
rect 10148 13028 10152 13084
rect 10088 13024 10152 13028
rect 14296 13084 14360 13088
rect 14296 13028 14300 13084
rect 14300 13028 14356 13084
rect 14356 13028 14360 13084
rect 14296 13024 14360 13028
rect 14376 13084 14440 13088
rect 14376 13028 14380 13084
rect 14380 13028 14436 13084
rect 14436 13028 14440 13084
rect 14376 13024 14440 13028
rect 14456 13084 14520 13088
rect 14456 13028 14460 13084
rect 14460 13028 14516 13084
rect 14516 13028 14520 13084
rect 14456 13024 14520 13028
rect 14536 13084 14600 13088
rect 14536 13028 14540 13084
rect 14540 13028 14596 13084
rect 14596 13028 14600 13084
rect 14536 13024 14600 13028
rect 3176 12540 3240 12544
rect 3176 12484 3180 12540
rect 3180 12484 3236 12540
rect 3236 12484 3240 12540
rect 3176 12480 3240 12484
rect 3256 12540 3320 12544
rect 3256 12484 3260 12540
rect 3260 12484 3316 12540
rect 3316 12484 3320 12540
rect 3256 12480 3320 12484
rect 3336 12540 3400 12544
rect 3336 12484 3340 12540
rect 3340 12484 3396 12540
rect 3396 12484 3400 12540
rect 3336 12480 3400 12484
rect 3416 12540 3480 12544
rect 3416 12484 3420 12540
rect 3420 12484 3476 12540
rect 3476 12484 3480 12540
rect 3416 12480 3480 12484
rect 7624 12540 7688 12544
rect 7624 12484 7628 12540
rect 7628 12484 7684 12540
rect 7684 12484 7688 12540
rect 7624 12480 7688 12484
rect 7704 12540 7768 12544
rect 7704 12484 7708 12540
rect 7708 12484 7764 12540
rect 7764 12484 7768 12540
rect 7704 12480 7768 12484
rect 7784 12540 7848 12544
rect 7784 12484 7788 12540
rect 7788 12484 7844 12540
rect 7844 12484 7848 12540
rect 7784 12480 7848 12484
rect 7864 12540 7928 12544
rect 7864 12484 7868 12540
rect 7868 12484 7924 12540
rect 7924 12484 7928 12540
rect 7864 12480 7928 12484
rect 12072 12540 12136 12544
rect 12072 12484 12076 12540
rect 12076 12484 12132 12540
rect 12132 12484 12136 12540
rect 12072 12480 12136 12484
rect 12152 12540 12216 12544
rect 12152 12484 12156 12540
rect 12156 12484 12212 12540
rect 12212 12484 12216 12540
rect 12152 12480 12216 12484
rect 12232 12540 12296 12544
rect 12232 12484 12236 12540
rect 12236 12484 12292 12540
rect 12292 12484 12296 12540
rect 12232 12480 12296 12484
rect 12312 12540 12376 12544
rect 12312 12484 12316 12540
rect 12316 12484 12372 12540
rect 12372 12484 12376 12540
rect 12312 12480 12376 12484
rect 16520 12540 16584 12544
rect 16520 12484 16524 12540
rect 16524 12484 16580 12540
rect 16580 12484 16584 12540
rect 16520 12480 16584 12484
rect 16600 12540 16664 12544
rect 16600 12484 16604 12540
rect 16604 12484 16660 12540
rect 16660 12484 16664 12540
rect 16600 12480 16664 12484
rect 16680 12540 16744 12544
rect 16680 12484 16684 12540
rect 16684 12484 16740 12540
rect 16740 12484 16744 12540
rect 16680 12480 16744 12484
rect 16760 12540 16824 12544
rect 16760 12484 16764 12540
rect 16764 12484 16820 12540
rect 16820 12484 16824 12540
rect 16760 12480 16824 12484
rect 5400 11996 5464 12000
rect 5400 11940 5404 11996
rect 5404 11940 5460 11996
rect 5460 11940 5464 11996
rect 5400 11936 5464 11940
rect 5480 11996 5544 12000
rect 5480 11940 5484 11996
rect 5484 11940 5540 11996
rect 5540 11940 5544 11996
rect 5480 11936 5544 11940
rect 5560 11996 5624 12000
rect 5560 11940 5564 11996
rect 5564 11940 5620 11996
rect 5620 11940 5624 11996
rect 5560 11936 5624 11940
rect 5640 11996 5704 12000
rect 5640 11940 5644 11996
rect 5644 11940 5700 11996
rect 5700 11940 5704 11996
rect 5640 11936 5704 11940
rect 9848 11996 9912 12000
rect 9848 11940 9852 11996
rect 9852 11940 9908 11996
rect 9908 11940 9912 11996
rect 9848 11936 9912 11940
rect 9928 11996 9992 12000
rect 9928 11940 9932 11996
rect 9932 11940 9988 11996
rect 9988 11940 9992 11996
rect 9928 11936 9992 11940
rect 10008 11996 10072 12000
rect 10008 11940 10012 11996
rect 10012 11940 10068 11996
rect 10068 11940 10072 11996
rect 10008 11936 10072 11940
rect 10088 11996 10152 12000
rect 10088 11940 10092 11996
rect 10092 11940 10148 11996
rect 10148 11940 10152 11996
rect 10088 11936 10152 11940
rect 14296 11996 14360 12000
rect 14296 11940 14300 11996
rect 14300 11940 14356 11996
rect 14356 11940 14360 11996
rect 14296 11936 14360 11940
rect 14376 11996 14440 12000
rect 14376 11940 14380 11996
rect 14380 11940 14436 11996
rect 14436 11940 14440 11996
rect 14376 11936 14440 11940
rect 14456 11996 14520 12000
rect 14456 11940 14460 11996
rect 14460 11940 14516 11996
rect 14516 11940 14520 11996
rect 14456 11936 14520 11940
rect 14536 11996 14600 12000
rect 14536 11940 14540 11996
rect 14540 11940 14596 11996
rect 14596 11940 14600 11996
rect 14536 11936 14600 11940
rect 3176 11452 3240 11456
rect 3176 11396 3180 11452
rect 3180 11396 3236 11452
rect 3236 11396 3240 11452
rect 3176 11392 3240 11396
rect 3256 11452 3320 11456
rect 3256 11396 3260 11452
rect 3260 11396 3316 11452
rect 3316 11396 3320 11452
rect 3256 11392 3320 11396
rect 3336 11452 3400 11456
rect 3336 11396 3340 11452
rect 3340 11396 3396 11452
rect 3396 11396 3400 11452
rect 3336 11392 3400 11396
rect 3416 11452 3480 11456
rect 3416 11396 3420 11452
rect 3420 11396 3476 11452
rect 3476 11396 3480 11452
rect 3416 11392 3480 11396
rect 7624 11452 7688 11456
rect 7624 11396 7628 11452
rect 7628 11396 7684 11452
rect 7684 11396 7688 11452
rect 7624 11392 7688 11396
rect 7704 11452 7768 11456
rect 7704 11396 7708 11452
rect 7708 11396 7764 11452
rect 7764 11396 7768 11452
rect 7704 11392 7768 11396
rect 7784 11452 7848 11456
rect 7784 11396 7788 11452
rect 7788 11396 7844 11452
rect 7844 11396 7848 11452
rect 7784 11392 7848 11396
rect 7864 11452 7928 11456
rect 7864 11396 7868 11452
rect 7868 11396 7924 11452
rect 7924 11396 7928 11452
rect 7864 11392 7928 11396
rect 12072 11452 12136 11456
rect 12072 11396 12076 11452
rect 12076 11396 12132 11452
rect 12132 11396 12136 11452
rect 12072 11392 12136 11396
rect 12152 11452 12216 11456
rect 12152 11396 12156 11452
rect 12156 11396 12212 11452
rect 12212 11396 12216 11452
rect 12152 11392 12216 11396
rect 12232 11452 12296 11456
rect 12232 11396 12236 11452
rect 12236 11396 12292 11452
rect 12292 11396 12296 11452
rect 12232 11392 12296 11396
rect 12312 11452 12376 11456
rect 12312 11396 12316 11452
rect 12316 11396 12372 11452
rect 12372 11396 12376 11452
rect 12312 11392 12376 11396
rect 16520 11452 16584 11456
rect 16520 11396 16524 11452
rect 16524 11396 16580 11452
rect 16580 11396 16584 11452
rect 16520 11392 16584 11396
rect 16600 11452 16664 11456
rect 16600 11396 16604 11452
rect 16604 11396 16660 11452
rect 16660 11396 16664 11452
rect 16600 11392 16664 11396
rect 16680 11452 16744 11456
rect 16680 11396 16684 11452
rect 16684 11396 16740 11452
rect 16740 11396 16744 11452
rect 16680 11392 16744 11396
rect 16760 11452 16824 11456
rect 16760 11396 16764 11452
rect 16764 11396 16820 11452
rect 16820 11396 16824 11452
rect 16760 11392 16824 11396
rect 5400 10908 5464 10912
rect 5400 10852 5404 10908
rect 5404 10852 5460 10908
rect 5460 10852 5464 10908
rect 5400 10848 5464 10852
rect 5480 10908 5544 10912
rect 5480 10852 5484 10908
rect 5484 10852 5540 10908
rect 5540 10852 5544 10908
rect 5480 10848 5544 10852
rect 5560 10908 5624 10912
rect 5560 10852 5564 10908
rect 5564 10852 5620 10908
rect 5620 10852 5624 10908
rect 5560 10848 5624 10852
rect 5640 10908 5704 10912
rect 5640 10852 5644 10908
rect 5644 10852 5700 10908
rect 5700 10852 5704 10908
rect 5640 10848 5704 10852
rect 9848 10908 9912 10912
rect 9848 10852 9852 10908
rect 9852 10852 9908 10908
rect 9908 10852 9912 10908
rect 9848 10848 9912 10852
rect 9928 10908 9992 10912
rect 9928 10852 9932 10908
rect 9932 10852 9988 10908
rect 9988 10852 9992 10908
rect 9928 10848 9992 10852
rect 10008 10908 10072 10912
rect 10008 10852 10012 10908
rect 10012 10852 10068 10908
rect 10068 10852 10072 10908
rect 10008 10848 10072 10852
rect 10088 10908 10152 10912
rect 10088 10852 10092 10908
rect 10092 10852 10148 10908
rect 10148 10852 10152 10908
rect 10088 10848 10152 10852
rect 14296 10908 14360 10912
rect 14296 10852 14300 10908
rect 14300 10852 14356 10908
rect 14356 10852 14360 10908
rect 14296 10848 14360 10852
rect 14376 10908 14440 10912
rect 14376 10852 14380 10908
rect 14380 10852 14436 10908
rect 14436 10852 14440 10908
rect 14376 10848 14440 10852
rect 14456 10908 14520 10912
rect 14456 10852 14460 10908
rect 14460 10852 14516 10908
rect 14516 10852 14520 10908
rect 14456 10848 14520 10852
rect 14536 10908 14600 10912
rect 14536 10852 14540 10908
rect 14540 10852 14596 10908
rect 14596 10852 14600 10908
rect 14536 10848 14600 10852
rect 3176 10364 3240 10368
rect 3176 10308 3180 10364
rect 3180 10308 3236 10364
rect 3236 10308 3240 10364
rect 3176 10304 3240 10308
rect 3256 10364 3320 10368
rect 3256 10308 3260 10364
rect 3260 10308 3316 10364
rect 3316 10308 3320 10364
rect 3256 10304 3320 10308
rect 3336 10364 3400 10368
rect 3336 10308 3340 10364
rect 3340 10308 3396 10364
rect 3396 10308 3400 10364
rect 3336 10304 3400 10308
rect 3416 10364 3480 10368
rect 3416 10308 3420 10364
rect 3420 10308 3476 10364
rect 3476 10308 3480 10364
rect 3416 10304 3480 10308
rect 7624 10364 7688 10368
rect 7624 10308 7628 10364
rect 7628 10308 7684 10364
rect 7684 10308 7688 10364
rect 7624 10304 7688 10308
rect 7704 10364 7768 10368
rect 7704 10308 7708 10364
rect 7708 10308 7764 10364
rect 7764 10308 7768 10364
rect 7704 10304 7768 10308
rect 7784 10364 7848 10368
rect 7784 10308 7788 10364
rect 7788 10308 7844 10364
rect 7844 10308 7848 10364
rect 7784 10304 7848 10308
rect 7864 10364 7928 10368
rect 7864 10308 7868 10364
rect 7868 10308 7924 10364
rect 7924 10308 7928 10364
rect 7864 10304 7928 10308
rect 12072 10364 12136 10368
rect 12072 10308 12076 10364
rect 12076 10308 12132 10364
rect 12132 10308 12136 10364
rect 12072 10304 12136 10308
rect 12152 10364 12216 10368
rect 12152 10308 12156 10364
rect 12156 10308 12212 10364
rect 12212 10308 12216 10364
rect 12152 10304 12216 10308
rect 12232 10364 12296 10368
rect 12232 10308 12236 10364
rect 12236 10308 12292 10364
rect 12292 10308 12296 10364
rect 12232 10304 12296 10308
rect 12312 10364 12376 10368
rect 12312 10308 12316 10364
rect 12316 10308 12372 10364
rect 12372 10308 12376 10364
rect 12312 10304 12376 10308
rect 16520 10364 16584 10368
rect 16520 10308 16524 10364
rect 16524 10308 16580 10364
rect 16580 10308 16584 10364
rect 16520 10304 16584 10308
rect 16600 10364 16664 10368
rect 16600 10308 16604 10364
rect 16604 10308 16660 10364
rect 16660 10308 16664 10364
rect 16600 10304 16664 10308
rect 16680 10364 16744 10368
rect 16680 10308 16684 10364
rect 16684 10308 16740 10364
rect 16740 10308 16744 10364
rect 16680 10304 16744 10308
rect 16760 10364 16824 10368
rect 16760 10308 16764 10364
rect 16764 10308 16820 10364
rect 16820 10308 16824 10364
rect 16760 10304 16824 10308
rect 5400 9820 5464 9824
rect 5400 9764 5404 9820
rect 5404 9764 5460 9820
rect 5460 9764 5464 9820
rect 5400 9760 5464 9764
rect 5480 9820 5544 9824
rect 5480 9764 5484 9820
rect 5484 9764 5540 9820
rect 5540 9764 5544 9820
rect 5480 9760 5544 9764
rect 5560 9820 5624 9824
rect 5560 9764 5564 9820
rect 5564 9764 5620 9820
rect 5620 9764 5624 9820
rect 5560 9760 5624 9764
rect 5640 9820 5704 9824
rect 5640 9764 5644 9820
rect 5644 9764 5700 9820
rect 5700 9764 5704 9820
rect 5640 9760 5704 9764
rect 9848 9820 9912 9824
rect 9848 9764 9852 9820
rect 9852 9764 9908 9820
rect 9908 9764 9912 9820
rect 9848 9760 9912 9764
rect 9928 9820 9992 9824
rect 9928 9764 9932 9820
rect 9932 9764 9988 9820
rect 9988 9764 9992 9820
rect 9928 9760 9992 9764
rect 10008 9820 10072 9824
rect 10008 9764 10012 9820
rect 10012 9764 10068 9820
rect 10068 9764 10072 9820
rect 10008 9760 10072 9764
rect 10088 9820 10152 9824
rect 10088 9764 10092 9820
rect 10092 9764 10148 9820
rect 10148 9764 10152 9820
rect 10088 9760 10152 9764
rect 14296 9820 14360 9824
rect 14296 9764 14300 9820
rect 14300 9764 14356 9820
rect 14356 9764 14360 9820
rect 14296 9760 14360 9764
rect 14376 9820 14440 9824
rect 14376 9764 14380 9820
rect 14380 9764 14436 9820
rect 14436 9764 14440 9820
rect 14376 9760 14440 9764
rect 14456 9820 14520 9824
rect 14456 9764 14460 9820
rect 14460 9764 14516 9820
rect 14516 9764 14520 9820
rect 14456 9760 14520 9764
rect 14536 9820 14600 9824
rect 14536 9764 14540 9820
rect 14540 9764 14596 9820
rect 14596 9764 14600 9820
rect 14536 9760 14600 9764
rect 3176 9276 3240 9280
rect 3176 9220 3180 9276
rect 3180 9220 3236 9276
rect 3236 9220 3240 9276
rect 3176 9216 3240 9220
rect 3256 9276 3320 9280
rect 3256 9220 3260 9276
rect 3260 9220 3316 9276
rect 3316 9220 3320 9276
rect 3256 9216 3320 9220
rect 3336 9276 3400 9280
rect 3336 9220 3340 9276
rect 3340 9220 3396 9276
rect 3396 9220 3400 9276
rect 3336 9216 3400 9220
rect 3416 9276 3480 9280
rect 3416 9220 3420 9276
rect 3420 9220 3476 9276
rect 3476 9220 3480 9276
rect 3416 9216 3480 9220
rect 7624 9276 7688 9280
rect 7624 9220 7628 9276
rect 7628 9220 7684 9276
rect 7684 9220 7688 9276
rect 7624 9216 7688 9220
rect 7704 9276 7768 9280
rect 7704 9220 7708 9276
rect 7708 9220 7764 9276
rect 7764 9220 7768 9276
rect 7704 9216 7768 9220
rect 7784 9276 7848 9280
rect 7784 9220 7788 9276
rect 7788 9220 7844 9276
rect 7844 9220 7848 9276
rect 7784 9216 7848 9220
rect 7864 9276 7928 9280
rect 7864 9220 7868 9276
rect 7868 9220 7924 9276
rect 7924 9220 7928 9276
rect 7864 9216 7928 9220
rect 12072 9276 12136 9280
rect 12072 9220 12076 9276
rect 12076 9220 12132 9276
rect 12132 9220 12136 9276
rect 12072 9216 12136 9220
rect 12152 9276 12216 9280
rect 12152 9220 12156 9276
rect 12156 9220 12212 9276
rect 12212 9220 12216 9276
rect 12152 9216 12216 9220
rect 12232 9276 12296 9280
rect 12232 9220 12236 9276
rect 12236 9220 12292 9276
rect 12292 9220 12296 9276
rect 12232 9216 12296 9220
rect 12312 9276 12376 9280
rect 12312 9220 12316 9276
rect 12316 9220 12372 9276
rect 12372 9220 12376 9276
rect 12312 9216 12376 9220
rect 16520 9276 16584 9280
rect 16520 9220 16524 9276
rect 16524 9220 16580 9276
rect 16580 9220 16584 9276
rect 16520 9216 16584 9220
rect 16600 9276 16664 9280
rect 16600 9220 16604 9276
rect 16604 9220 16660 9276
rect 16660 9220 16664 9276
rect 16600 9216 16664 9220
rect 16680 9276 16744 9280
rect 16680 9220 16684 9276
rect 16684 9220 16740 9276
rect 16740 9220 16744 9276
rect 16680 9216 16744 9220
rect 16760 9276 16824 9280
rect 16760 9220 16764 9276
rect 16764 9220 16820 9276
rect 16820 9220 16824 9276
rect 16760 9216 16824 9220
rect 5400 8732 5464 8736
rect 5400 8676 5404 8732
rect 5404 8676 5460 8732
rect 5460 8676 5464 8732
rect 5400 8672 5464 8676
rect 5480 8732 5544 8736
rect 5480 8676 5484 8732
rect 5484 8676 5540 8732
rect 5540 8676 5544 8732
rect 5480 8672 5544 8676
rect 5560 8732 5624 8736
rect 5560 8676 5564 8732
rect 5564 8676 5620 8732
rect 5620 8676 5624 8732
rect 5560 8672 5624 8676
rect 5640 8732 5704 8736
rect 5640 8676 5644 8732
rect 5644 8676 5700 8732
rect 5700 8676 5704 8732
rect 5640 8672 5704 8676
rect 9848 8732 9912 8736
rect 9848 8676 9852 8732
rect 9852 8676 9908 8732
rect 9908 8676 9912 8732
rect 9848 8672 9912 8676
rect 9928 8732 9992 8736
rect 9928 8676 9932 8732
rect 9932 8676 9988 8732
rect 9988 8676 9992 8732
rect 9928 8672 9992 8676
rect 10008 8732 10072 8736
rect 10008 8676 10012 8732
rect 10012 8676 10068 8732
rect 10068 8676 10072 8732
rect 10008 8672 10072 8676
rect 10088 8732 10152 8736
rect 10088 8676 10092 8732
rect 10092 8676 10148 8732
rect 10148 8676 10152 8732
rect 10088 8672 10152 8676
rect 14296 8732 14360 8736
rect 14296 8676 14300 8732
rect 14300 8676 14356 8732
rect 14356 8676 14360 8732
rect 14296 8672 14360 8676
rect 14376 8732 14440 8736
rect 14376 8676 14380 8732
rect 14380 8676 14436 8732
rect 14436 8676 14440 8732
rect 14376 8672 14440 8676
rect 14456 8732 14520 8736
rect 14456 8676 14460 8732
rect 14460 8676 14516 8732
rect 14516 8676 14520 8732
rect 14456 8672 14520 8676
rect 14536 8732 14600 8736
rect 14536 8676 14540 8732
rect 14540 8676 14596 8732
rect 14596 8676 14600 8732
rect 14536 8672 14600 8676
rect 3176 8188 3240 8192
rect 3176 8132 3180 8188
rect 3180 8132 3236 8188
rect 3236 8132 3240 8188
rect 3176 8128 3240 8132
rect 3256 8188 3320 8192
rect 3256 8132 3260 8188
rect 3260 8132 3316 8188
rect 3316 8132 3320 8188
rect 3256 8128 3320 8132
rect 3336 8188 3400 8192
rect 3336 8132 3340 8188
rect 3340 8132 3396 8188
rect 3396 8132 3400 8188
rect 3336 8128 3400 8132
rect 3416 8188 3480 8192
rect 3416 8132 3420 8188
rect 3420 8132 3476 8188
rect 3476 8132 3480 8188
rect 3416 8128 3480 8132
rect 7624 8188 7688 8192
rect 7624 8132 7628 8188
rect 7628 8132 7684 8188
rect 7684 8132 7688 8188
rect 7624 8128 7688 8132
rect 7704 8188 7768 8192
rect 7704 8132 7708 8188
rect 7708 8132 7764 8188
rect 7764 8132 7768 8188
rect 7704 8128 7768 8132
rect 7784 8188 7848 8192
rect 7784 8132 7788 8188
rect 7788 8132 7844 8188
rect 7844 8132 7848 8188
rect 7784 8128 7848 8132
rect 7864 8188 7928 8192
rect 7864 8132 7868 8188
rect 7868 8132 7924 8188
rect 7924 8132 7928 8188
rect 7864 8128 7928 8132
rect 12072 8188 12136 8192
rect 12072 8132 12076 8188
rect 12076 8132 12132 8188
rect 12132 8132 12136 8188
rect 12072 8128 12136 8132
rect 12152 8188 12216 8192
rect 12152 8132 12156 8188
rect 12156 8132 12212 8188
rect 12212 8132 12216 8188
rect 12152 8128 12216 8132
rect 12232 8188 12296 8192
rect 12232 8132 12236 8188
rect 12236 8132 12292 8188
rect 12292 8132 12296 8188
rect 12232 8128 12296 8132
rect 12312 8188 12376 8192
rect 12312 8132 12316 8188
rect 12316 8132 12372 8188
rect 12372 8132 12376 8188
rect 12312 8128 12376 8132
rect 16520 8188 16584 8192
rect 16520 8132 16524 8188
rect 16524 8132 16580 8188
rect 16580 8132 16584 8188
rect 16520 8128 16584 8132
rect 16600 8188 16664 8192
rect 16600 8132 16604 8188
rect 16604 8132 16660 8188
rect 16660 8132 16664 8188
rect 16600 8128 16664 8132
rect 16680 8188 16744 8192
rect 16680 8132 16684 8188
rect 16684 8132 16740 8188
rect 16740 8132 16744 8188
rect 16680 8128 16744 8132
rect 16760 8188 16824 8192
rect 16760 8132 16764 8188
rect 16764 8132 16820 8188
rect 16820 8132 16824 8188
rect 16760 8128 16824 8132
rect 5400 7644 5464 7648
rect 5400 7588 5404 7644
rect 5404 7588 5460 7644
rect 5460 7588 5464 7644
rect 5400 7584 5464 7588
rect 5480 7644 5544 7648
rect 5480 7588 5484 7644
rect 5484 7588 5540 7644
rect 5540 7588 5544 7644
rect 5480 7584 5544 7588
rect 5560 7644 5624 7648
rect 5560 7588 5564 7644
rect 5564 7588 5620 7644
rect 5620 7588 5624 7644
rect 5560 7584 5624 7588
rect 5640 7644 5704 7648
rect 5640 7588 5644 7644
rect 5644 7588 5700 7644
rect 5700 7588 5704 7644
rect 5640 7584 5704 7588
rect 9848 7644 9912 7648
rect 9848 7588 9852 7644
rect 9852 7588 9908 7644
rect 9908 7588 9912 7644
rect 9848 7584 9912 7588
rect 9928 7644 9992 7648
rect 9928 7588 9932 7644
rect 9932 7588 9988 7644
rect 9988 7588 9992 7644
rect 9928 7584 9992 7588
rect 10008 7644 10072 7648
rect 10008 7588 10012 7644
rect 10012 7588 10068 7644
rect 10068 7588 10072 7644
rect 10008 7584 10072 7588
rect 10088 7644 10152 7648
rect 10088 7588 10092 7644
rect 10092 7588 10148 7644
rect 10148 7588 10152 7644
rect 10088 7584 10152 7588
rect 14296 7644 14360 7648
rect 14296 7588 14300 7644
rect 14300 7588 14356 7644
rect 14356 7588 14360 7644
rect 14296 7584 14360 7588
rect 14376 7644 14440 7648
rect 14376 7588 14380 7644
rect 14380 7588 14436 7644
rect 14436 7588 14440 7644
rect 14376 7584 14440 7588
rect 14456 7644 14520 7648
rect 14456 7588 14460 7644
rect 14460 7588 14516 7644
rect 14516 7588 14520 7644
rect 14456 7584 14520 7588
rect 14536 7644 14600 7648
rect 14536 7588 14540 7644
rect 14540 7588 14596 7644
rect 14596 7588 14600 7644
rect 14536 7584 14600 7588
rect 3176 7100 3240 7104
rect 3176 7044 3180 7100
rect 3180 7044 3236 7100
rect 3236 7044 3240 7100
rect 3176 7040 3240 7044
rect 3256 7100 3320 7104
rect 3256 7044 3260 7100
rect 3260 7044 3316 7100
rect 3316 7044 3320 7100
rect 3256 7040 3320 7044
rect 3336 7100 3400 7104
rect 3336 7044 3340 7100
rect 3340 7044 3396 7100
rect 3396 7044 3400 7100
rect 3336 7040 3400 7044
rect 3416 7100 3480 7104
rect 3416 7044 3420 7100
rect 3420 7044 3476 7100
rect 3476 7044 3480 7100
rect 3416 7040 3480 7044
rect 7624 7100 7688 7104
rect 7624 7044 7628 7100
rect 7628 7044 7684 7100
rect 7684 7044 7688 7100
rect 7624 7040 7688 7044
rect 7704 7100 7768 7104
rect 7704 7044 7708 7100
rect 7708 7044 7764 7100
rect 7764 7044 7768 7100
rect 7704 7040 7768 7044
rect 7784 7100 7848 7104
rect 7784 7044 7788 7100
rect 7788 7044 7844 7100
rect 7844 7044 7848 7100
rect 7784 7040 7848 7044
rect 7864 7100 7928 7104
rect 7864 7044 7868 7100
rect 7868 7044 7924 7100
rect 7924 7044 7928 7100
rect 7864 7040 7928 7044
rect 12072 7100 12136 7104
rect 12072 7044 12076 7100
rect 12076 7044 12132 7100
rect 12132 7044 12136 7100
rect 12072 7040 12136 7044
rect 12152 7100 12216 7104
rect 12152 7044 12156 7100
rect 12156 7044 12212 7100
rect 12212 7044 12216 7100
rect 12152 7040 12216 7044
rect 12232 7100 12296 7104
rect 12232 7044 12236 7100
rect 12236 7044 12292 7100
rect 12292 7044 12296 7100
rect 12232 7040 12296 7044
rect 12312 7100 12376 7104
rect 12312 7044 12316 7100
rect 12316 7044 12372 7100
rect 12372 7044 12376 7100
rect 12312 7040 12376 7044
rect 16520 7100 16584 7104
rect 16520 7044 16524 7100
rect 16524 7044 16580 7100
rect 16580 7044 16584 7100
rect 16520 7040 16584 7044
rect 16600 7100 16664 7104
rect 16600 7044 16604 7100
rect 16604 7044 16660 7100
rect 16660 7044 16664 7100
rect 16600 7040 16664 7044
rect 16680 7100 16744 7104
rect 16680 7044 16684 7100
rect 16684 7044 16740 7100
rect 16740 7044 16744 7100
rect 16680 7040 16744 7044
rect 16760 7100 16824 7104
rect 16760 7044 16764 7100
rect 16764 7044 16820 7100
rect 16820 7044 16824 7100
rect 16760 7040 16824 7044
rect 5400 6556 5464 6560
rect 5400 6500 5404 6556
rect 5404 6500 5460 6556
rect 5460 6500 5464 6556
rect 5400 6496 5464 6500
rect 5480 6556 5544 6560
rect 5480 6500 5484 6556
rect 5484 6500 5540 6556
rect 5540 6500 5544 6556
rect 5480 6496 5544 6500
rect 5560 6556 5624 6560
rect 5560 6500 5564 6556
rect 5564 6500 5620 6556
rect 5620 6500 5624 6556
rect 5560 6496 5624 6500
rect 5640 6556 5704 6560
rect 5640 6500 5644 6556
rect 5644 6500 5700 6556
rect 5700 6500 5704 6556
rect 5640 6496 5704 6500
rect 9848 6556 9912 6560
rect 9848 6500 9852 6556
rect 9852 6500 9908 6556
rect 9908 6500 9912 6556
rect 9848 6496 9912 6500
rect 9928 6556 9992 6560
rect 9928 6500 9932 6556
rect 9932 6500 9988 6556
rect 9988 6500 9992 6556
rect 9928 6496 9992 6500
rect 10008 6556 10072 6560
rect 10008 6500 10012 6556
rect 10012 6500 10068 6556
rect 10068 6500 10072 6556
rect 10008 6496 10072 6500
rect 10088 6556 10152 6560
rect 10088 6500 10092 6556
rect 10092 6500 10148 6556
rect 10148 6500 10152 6556
rect 10088 6496 10152 6500
rect 14296 6556 14360 6560
rect 14296 6500 14300 6556
rect 14300 6500 14356 6556
rect 14356 6500 14360 6556
rect 14296 6496 14360 6500
rect 14376 6556 14440 6560
rect 14376 6500 14380 6556
rect 14380 6500 14436 6556
rect 14436 6500 14440 6556
rect 14376 6496 14440 6500
rect 14456 6556 14520 6560
rect 14456 6500 14460 6556
rect 14460 6500 14516 6556
rect 14516 6500 14520 6556
rect 14456 6496 14520 6500
rect 14536 6556 14600 6560
rect 14536 6500 14540 6556
rect 14540 6500 14596 6556
rect 14596 6500 14600 6556
rect 14536 6496 14600 6500
rect 3176 6012 3240 6016
rect 3176 5956 3180 6012
rect 3180 5956 3236 6012
rect 3236 5956 3240 6012
rect 3176 5952 3240 5956
rect 3256 6012 3320 6016
rect 3256 5956 3260 6012
rect 3260 5956 3316 6012
rect 3316 5956 3320 6012
rect 3256 5952 3320 5956
rect 3336 6012 3400 6016
rect 3336 5956 3340 6012
rect 3340 5956 3396 6012
rect 3396 5956 3400 6012
rect 3336 5952 3400 5956
rect 3416 6012 3480 6016
rect 3416 5956 3420 6012
rect 3420 5956 3476 6012
rect 3476 5956 3480 6012
rect 3416 5952 3480 5956
rect 7624 6012 7688 6016
rect 7624 5956 7628 6012
rect 7628 5956 7684 6012
rect 7684 5956 7688 6012
rect 7624 5952 7688 5956
rect 7704 6012 7768 6016
rect 7704 5956 7708 6012
rect 7708 5956 7764 6012
rect 7764 5956 7768 6012
rect 7704 5952 7768 5956
rect 7784 6012 7848 6016
rect 7784 5956 7788 6012
rect 7788 5956 7844 6012
rect 7844 5956 7848 6012
rect 7784 5952 7848 5956
rect 7864 6012 7928 6016
rect 7864 5956 7868 6012
rect 7868 5956 7924 6012
rect 7924 5956 7928 6012
rect 7864 5952 7928 5956
rect 12072 6012 12136 6016
rect 12072 5956 12076 6012
rect 12076 5956 12132 6012
rect 12132 5956 12136 6012
rect 12072 5952 12136 5956
rect 12152 6012 12216 6016
rect 12152 5956 12156 6012
rect 12156 5956 12212 6012
rect 12212 5956 12216 6012
rect 12152 5952 12216 5956
rect 12232 6012 12296 6016
rect 12232 5956 12236 6012
rect 12236 5956 12292 6012
rect 12292 5956 12296 6012
rect 12232 5952 12296 5956
rect 12312 6012 12376 6016
rect 12312 5956 12316 6012
rect 12316 5956 12372 6012
rect 12372 5956 12376 6012
rect 12312 5952 12376 5956
rect 16520 6012 16584 6016
rect 16520 5956 16524 6012
rect 16524 5956 16580 6012
rect 16580 5956 16584 6012
rect 16520 5952 16584 5956
rect 16600 6012 16664 6016
rect 16600 5956 16604 6012
rect 16604 5956 16660 6012
rect 16660 5956 16664 6012
rect 16600 5952 16664 5956
rect 16680 6012 16744 6016
rect 16680 5956 16684 6012
rect 16684 5956 16740 6012
rect 16740 5956 16744 6012
rect 16680 5952 16744 5956
rect 16760 6012 16824 6016
rect 16760 5956 16764 6012
rect 16764 5956 16820 6012
rect 16820 5956 16824 6012
rect 16760 5952 16824 5956
rect 5400 5468 5464 5472
rect 5400 5412 5404 5468
rect 5404 5412 5460 5468
rect 5460 5412 5464 5468
rect 5400 5408 5464 5412
rect 5480 5468 5544 5472
rect 5480 5412 5484 5468
rect 5484 5412 5540 5468
rect 5540 5412 5544 5468
rect 5480 5408 5544 5412
rect 5560 5468 5624 5472
rect 5560 5412 5564 5468
rect 5564 5412 5620 5468
rect 5620 5412 5624 5468
rect 5560 5408 5624 5412
rect 5640 5468 5704 5472
rect 5640 5412 5644 5468
rect 5644 5412 5700 5468
rect 5700 5412 5704 5468
rect 5640 5408 5704 5412
rect 9848 5468 9912 5472
rect 9848 5412 9852 5468
rect 9852 5412 9908 5468
rect 9908 5412 9912 5468
rect 9848 5408 9912 5412
rect 9928 5468 9992 5472
rect 9928 5412 9932 5468
rect 9932 5412 9988 5468
rect 9988 5412 9992 5468
rect 9928 5408 9992 5412
rect 10008 5468 10072 5472
rect 10008 5412 10012 5468
rect 10012 5412 10068 5468
rect 10068 5412 10072 5468
rect 10008 5408 10072 5412
rect 10088 5468 10152 5472
rect 10088 5412 10092 5468
rect 10092 5412 10148 5468
rect 10148 5412 10152 5468
rect 10088 5408 10152 5412
rect 14296 5468 14360 5472
rect 14296 5412 14300 5468
rect 14300 5412 14356 5468
rect 14356 5412 14360 5468
rect 14296 5408 14360 5412
rect 14376 5468 14440 5472
rect 14376 5412 14380 5468
rect 14380 5412 14436 5468
rect 14436 5412 14440 5468
rect 14376 5408 14440 5412
rect 14456 5468 14520 5472
rect 14456 5412 14460 5468
rect 14460 5412 14516 5468
rect 14516 5412 14520 5468
rect 14456 5408 14520 5412
rect 14536 5468 14600 5472
rect 14536 5412 14540 5468
rect 14540 5412 14596 5468
rect 14596 5412 14600 5468
rect 14536 5408 14600 5412
rect 3176 4924 3240 4928
rect 3176 4868 3180 4924
rect 3180 4868 3236 4924
rect 3236 4868 3240 4924
rect 3176 4864 3240 4868
rect 3256 4924 3320 4928
rect 3256 4868 3260 4924
rect 3260 4868 3316 4924
rect 3316 4868 3320 4924
rect 3256 4864 3320 4868
rect 3336 4924 3400 4928
rect 3336 4868 3340 4924
rect 3340 4868 3396 4924
rect 3396 4868 3400 4924
rect 3336 4864 3400 4868
rect 3416 4924 3480 4928
rect 3416 4868 3420 4924
rect 3420 4868 3476 4924
rect 3476 4868 3480 4924
rect 3416 4864 3480 4868
rect 7624 4924 7688 4928
rect 7624 4868 7628 4924
rect 7628 4868 7684 4924
rect 7684 4868 7688 4924
rect 7624 4864 7688 4868
rect 7704 4924 7768 4928
rect 7704 4868 7708 4924
rect 7708 4868 7764 4924
rect 7764 4868 7768 4924
rect 7704 4864 7768 4868
rect 7784 4924 7848 4928
rect 7784 4868 7788 4924
rect 7788 4868 7844 4924
rect 7844 4868 7848 4924
rect 7784 4864 7848 4868
rect 7864 4924 7928 4928
rect 7864 4868 7868 4924
rect 7868 4868 7924 4924
rect 7924 4868 7928 4924
rect 7864 4864 7928 4868
rect 12072 4924 12136 4928
rect 12072 4868 12076 4924
rect 12076 4868 12132 4924
rect 12132 4868 12136 4924
rect 12072 4864 12136 4868
rect 12152 4924 12216 4928
rect 12152 4868 12156 4924
rect 12156 4868 12212 4924
rect 12212 4868 12216 4924
rect 12152 4864 12216 4868
rect 12232 4924 12296 4928
rect 12232 4868 12236 4924
rect 12236 4868 12292 4924
rect 12292 4868 12296 4924
rect 12232 4864 12296 4868
rect 12312 4924 12376 4928
rect 12312 4868 12316 4924
rect 12316 4868 12372 4924
rect 12372 4868 12376 4924
rect 12312 4864 12376 4868
rect 16520 4924 16584 4928
rect 16520 4868 16524 4924
rect 16524 4868 16580 4924
rect 16580 4868 16584 4924
rect 16520 4864 16584 4868
rect 16600 4924 16664 4928
rect 16600 4868 16604 4924
rect 16604 4868 16660 4924
rect 16660 4868 16664 4924
rect 16600 4864 16664 4868
rect 16680 4924 16744 4928
rect 16680 4868 16684 4924
rect 16684 4868 16740 4924
rect 16740 4868 16744 4924
rect 16680 4864 16744 4868
rect 16760 4924 16824 4928
rect 16760 4868 16764 4924
rect 16764 4868 16820 4924
rect 16820 4868 16824 4924
rect 16760 4864 16824 4868
rect 5400 4380 5464 4384
rect 5400 4324 5404 4380
rect 5404 4324 5460 4380
rect 5460 4324 5464 4380
rect 5400 4320 5464 4324
rect 5480 4380 5544 4384
rect 5480 4324 5484 4380
rect 5484 4324 5540 4380
rect 5540 4324 5544 4380
rect 5480 4320 5544 4324
rect 5560 4380 5624 4384
rect 5560 4324 5564 4380
rect 5564 4324 5620 4380
rect 5620 4324 5624 4380
rect 5560 4320 5624 4324
rect 5640 4380 5704 4384
rect 5640 4324 5644 4380
rect 5644 4324 5700 4380
rect 5700 4324 5704 4380
rect 5640 4320 5704 4324
rect 9848 4380 9912 4384
rect 9848 4324 9852 4380
rect 9852 4324 9908 4380
rect 9908 4324 9912 4380
rect 9848 4320 9912 4324
rect 9928 4380 9992 4384
rect 9928 4324 9932 4380
rect 9932 4324 9988 4380
rect 9988 4324 9992 4380
rect 9928 4320 9992 4324
rect 10008 4380 10072 4384
rect 10008 4324 10012 4380
rect 10012 4324 10068 4380
rect 10068 4324 10072 4380
rect 10008 4320 10072 4324
rect 10088 4380 10152 4384
rect 10088 4324 10092 4380
rect 10092 4324 10148 4380
rect 10148 4324 10152 4380
rect 10088 4320 10152 4324
rect 14296 4380 14360 4384
rect 14296 4324 14300 4380
rect 14300 4324 14356 4380
rect 14356 4324 14360 4380
rect 14296 4320 14360 4324
rect 14376 4380 14440 4384
rect 14376 4324 14380 4380
rect 14380 4324 14436 4380
rect 14436 4324 14440 4380
rect 14376 4320 14440 4324
rect 14456 4380 14520 4384
rect 14456 4324 14460 4380
rect 14460 4324 14516 4380
rect 14516 4324 14520 4380
rect 14456 4320 14520 4324
rect 14536 4380 14600 4384
rect 14536 4324 14540 4380
rect 14540 4324 14596 4380
rect 14596 4324 14600 4380
rect 14536 4320 14600 4324
rect 3176 3836 3240 3840
rect 3176 3780 3180 3836
rect 3180 3780 3236 3836
rect 3236 3780 3240 3836
rect 3176 3776 3240 3780
rect 3256 3836 3320 3840
rect 3256 3780 3260 3836
rect 3260 3780 3316 3836
rect 3316 3780 3320 3836
rect 3256 3776 3320 3780
rect 3336 3836 3400 3840
rect 3336 3780 3340 3836
rect 3340 3780 3396 3836
rect 3396 3780 3400 3836
rect 3336 3776 3400 3780
rect 3416 3836 3480 3840
rect 3416 3780 3420 3836
rect 3420 3780 3476 3836
rect 3476 3780 3480 3836
rect 3416 3776 3480 3780
rect 7624 3836 7688 3840
rect 7624 3780 7628 3836
rect 7628 3780 7684 3836
rect 7684 3780 7688 3836
rect 7624 3776 7688 3780
rect 7704 3836 7768 3840
rect 7704 3780 7708 3836
rect 7708 3780 7764 3836
rect 7764 3780 7768 3836
rect 7704 3776 7768 3780
rect 7784 3836 7848 3840
rect 7784 3780 7788 3836
rect 7788 3780 7844 3836
rect 7844 3780 7848 3836
rect 7784 3776 7848 3780
rect 7864 3836 7928 3840
rect 7864 3780 7868 3836
rect 7868 3780 7924 3836
rect 7924 3780 7928 3836
rect 7864 3776 7928 3780
rect 12072 3836 12136 3840
rect 12072 3780 12076 3836
rect 12076 3780 12132 3836
rect 12132 3780 12136 3836
rect 12072 3776 12136 3780
rect 12152 3836 12216 3840
rect 12152 3780 12156 3836
rect 12156 3780 12212 3836
rect 12212 3780 12216 3836
rect 12152 3776 12216 3780
rect 12232 3836 12296 3840
rect 12232 3780 12236 3836
rect 12236 3780 12292 3836
rect 12292 3780 12296 3836
rect 12232 3776 12296 3780
rect 12312 3836 12376 3840
rect 12312 3780 12316 3836
rect 12316 3780 12372 3836
rect 12372 3780 12376 3836
rect 12312 3776 12376 3780
rect 16520 3836 16584 3840
rect 16520 3780 16524 3836
rect 16524 3780 16580 3836
rect 16580 3780 16584 3836
rect 16520 3776 16584 3780
rect 16600 3836 16664 3840
rect 16600 3780 16604 3836
rect 16604 3780 16660 3836
rect 16660 3780 16664 3836
rect 16600 3776 16664 3780
rect 16680 3836 16744 3840
rect 16680 3780 16684 3836
rect 16684 3780 16740 3836
rect 16740 3780 16744 3836
rect 16680 3776 16744 3780
rect 16760 3836 16824 3840
rect 16760 3780 16764 3836
rect 16764 3780 16820 3836
rect 16820 3780 16824 3836
rect 16760 3776 16824 3780
rect 5400 3292 5464 3296
rect 5400 3236 5404 3292
rect 5404 3236 5460 3292
rect 5460 3236 5464 3292
rect 5400 3232 5464 3236
rect 5480 3292 5544 3296
rect 5480 3236 5484 3292
rect 5484 3236 5540 3292
rect 5540 3236 5544 3292
rect 5480 3232 5544 3236
rect 5560 3292 5624 3296
rect 5560 3236 5564 3292
rect 5564 3236 5620 3292
rect 5620 3236 5624 3292
rect 5560 3232 5624 3236
rect 5640 3292 5704 3296
rect 5640 3236 5644 3292
rect 5644 3236 5700 3292
rect 5700 3236 5704 3292
rect 5640 3232 5704 3236
rect 9848 3292 9912 3296
rect 9848 3236 9852 3292
rect 9852 3236 9908 3292
rect 9908 3236 9912 3292
rect 9848 3232 9912 3236
rect 9928 3292 9992 3296
rect 9928 3236 9932 3292
rect 9932 3236 9988 3292
rect 9988 3236 9992 3292
rect 9928 3232 9992 3236
rect 10008 3292 10072 3296
rect 10008 3236 10012 3292
rect 10012 3236 10068 3292
rect 10068 3236 10072 3292
rect 10008 3232 10072 3236
rect 10088 3292 10152 3296
rect 10088 3236 10092 3292
rect 10092 3236 10148 3292
rect 10148 3236 10152 3292
rect 10088 3232 10152 3236
rect 14296 3292 14360 3296
rect 14296 3236 14300 3292
rect 14300 3236 14356 3292
rect 14356 3236 14360 3292
rect 14296 3232 14360 3236
rect 14376 3292 14440 3296
rect 14376 3236 14380 3292
rect 14380 3236 14436 3292
rect 14436 3236 14440 3292
rect 14376 3232 14440 3236
rect 14456 3292 14520 3296
rect 14456 3236 14460 3292
rect 14460 3236 14516 3292
rect 14516 3236 14520 3292
rect 14456 3232 14520 3236
rect 14536 3292 14600 3296
rect 14536 3236 14540 3292
rect 14540 3236 14596 3292
rect 14596 3236 14600 3292
rect 14536 3232 14600 3236
rect 3176 2748 3240 2752
rect 3176 2692 3180 2748
rect 3180 2692 3236 2748
rect 3236 2692 3240 2748
rect 3176 2688 3240 2692
rect 3256 2748 3320 2752
rect 3256 2692 3260 2748
rect 3260 2692 3316 2748
rect 3316 2692 3320 2748
rect 3256 2688 3320 2692
rect 3336 2748 3400 2752
rect 3336 2692 3340 2748
rect 3340 2692 3396 2748
rect 3396 2692 3400 2748
rect 3336 2688 3400 2692
rect 3416 2748 3480 2752
rect 3416 2692 3420 2748
rect 3420 2692 3476 2748
rect 3476 2692 3480 2748
rect 3416 2688 3480 2692
rect 7624 2748 7688 2752
rect 7624 2692 7628 2748
rect 7628 2692 7684 2748
rect 7684 2692 7688 2748
rect 7624 2688 7688 2692
rect 7704 2748 7768 2752
rect 7704 2692 7708 2748
rect 7708 2692 7764 2748
rect 7764 2692 7768 2748
rect 7704 2688 7768 2692
rect 7784 2748 7848 2752
rect 7784 2692 7788 2748
rect 7788 2692 7844 2748
rect 7844 2692 7848 2748
rect 7784 2688 7848 2692
rect 7864 2748 7928 2752
rect 7864 2692 7868 2748
rect 7868 2692 7924 2748
rect 7924 2692 7928 2748
rect 7864 2688 7928 2692
rect 12072 2748 12136 2752
rect 12072 2692 12076 2748
rect 12076 2692 12132 2748
rect 12132 2692 12136 2748
rect 12072 2688 12136 2692
rect 12152 2748 12216 2752
rect 12152 2692 12156 2748
rect 12156 2692 12212 2748
rect 12212 2692 12216 2748
rect 12152 2688 12216 2692
rect 12232 2748 12296 2752
rect 12232 2692 12236 2748
rect 12236 2692 12292 2748
rect 12292 2692 12296 2748
rect 12232 2688 12296 2692
rect 12312 2748 12376 2752
rect 12312 2692 12316 2748
rect 12316 2692 12372 2748
rect 12372 2692 12376 2748
rect 12312 2688 12376 2692
rect 16520 2748 16584 2752
rect 16520 2692 16524 2748
rect 16524 2692 16580 2748
rect 16580 2692 16584 2748
rect 16520 2688 16584 2692
rect 16600 2748 16664 2752
rect 16600 2692 16604 2748
rect 16604 2692 16660 2748
rect 16660 2692 16664 2748
rect 16600 2688 16664 2692
rect 16680 2748 16744 2752
rect 16680 2692 16684 2748
rect 16684 2692 16740 2748
rect 16740 2692 16744 2748
rect 16680 2688 16744 2692
rect 16760 2748 16824 2752
rect 16760 2692 16764 2748
rect 16764 2692 16820 2748
rect 16820 2692 16824 2748
rect 16760 2688 16824 2692
rect 5400 2204 5464 2208
rect 5400 2148 5404 2204
rect 5404 2148 5460 2204
rect 5460 2148 5464 2204
rect 5400 2144 5464 2148
rect 5480 2204 5544 2208
rect 5480 2148 5484 2204
rect 5484 2148 5540 2204
rect 5540 2148 5544 2204
rect 5480 2144 5544 2148
rect 5560 2204 5624 2208
rect 5560 2148 5564 2204
rect 5564 2148 5620 2204
rect 5620 2148 5624 2204
rect 5560 2144 5624 2148
rect 5640 2204 5704 2208
rect 5640 2148 5644 2204
rect 5644 2148 5700 2204
rect 5700 2148 5704 2204
rect 5640 2144 5704 2148
rect 9848 2204 9912 2208
rect 9848 2148 9852 2204
rect 9852 2148 9908 2204
rect 9908 2148 9912 2204
rect 9848 2144 9912 2148
rect 9928 2204 9992 2208
rect 9928 2148 9932 2204
rect 9932 2148 9988 2204
rect 9988 2148 9992 2204
rect 9928 2144 9992 2148
rect 10008 2204 10072 2208
rect 10008 2148 10012 2204
rect 10012 2148 10068 2204
rect 10068 2148 10072 2204
rect 10008 2144 10072 2148
rect 10088 2204 10152 2208
rect 10088 2148 10092 2204
rect 10092 2148 10148 2204
rect 10148 2148 10152 2204
rect 10088 2144 10152 2148
rect 14296 2204 14360 2208
rect 14296 2148 14300 2204
rect 14300 2148 14356 2204
rect 14356 2148 14360 2204
rect 14296 2144 14360 2148
rect 14376 2204 14440 2208
rect 14376 2148 14380 2204
rect 14380 2148 14436 2204
rect 14436 2148 14440 2204
rect 14376 2144 14440 2148
rect 14456 2204 14520 2208
rect 14456 2148 14460 2204
rect 14460 2148 14516 2204
rect 14516 2148 14520 2204
rect 14456 2144 14520 2148
rect 14536 2204 14600 2208
rect 14536 2148 14540 2204
rect 14540 2148 14596 2204
rect 14596 2148 14600 2204
rect 14536 2144 14600 2148
<< metal4 >>
rect 3168 16896 3488 17456
rect 3168 16832 3176 16896
rect 3240 16832 3256 16896
rect 3320 16832 3336 16896
rect 3400 16832 3416 16896
rect 3480 16832 3488 16896
rect 3168 15986 3488 16832
rect 3168 15808 3210 15986
rect 3446 15808 3488 15986
rect 3168 15744 3176 15808
rect 3240 15744 3256 15750
rect 3320 15744 3336 15750
rect 3400 15744 3416 15750
rect 3480 15744 3488 15808
rect 3168 14720 3488 15744
rect 3168 14656 3176 14720
rect 3240 14656 3256 14720
rect 3320 14656 3336 14720
rect 3400 14656 3416 14720
rect 3480 14656 3488 14720
rect 3168 13632 3488 14656
rect 3168 13568 3176 13632
rect 3240 13568 3256 13632
rect 3320 13568 3336 13632
rect 3400 13568 3416 13632
rect 3480 13568 3488 13632
rect 3168 12544 3488 13568
rect 3168 12480 3176 12544
rect 3240 12480 3256 12544
rect 3320 12480 3336 12544
rect 3400 12480 3416 12544
rect 3480 12480 3488 12544
rect 3168 12074 3488 12480
rect 3168 11838 3210 12074
rect 3446 11838 3488 12074
rect 3168 11456 3488 11838
rect 3168 11392 3176 11456
rect 3240 11392 3256 11456
rect 3320 11392 3336 11456
rect 3400 11392 3416 11456
rect 3480 11392 3488 11456
rect 3168 10368 3488 11392
rect 3168 10304 3176 10368
rect 3240 10304 3256 10368
rect 3320 10304 3336 10368
rect 3400 10304 3416 10368
rect 3480 10304 3488 10368
rect 3168 9280 3488 10304
rect 3168 9216 3176 9280
rect 3240 9216 3256 9280
rect 3320 9216 3336 9280
rect 3400 9216 3416 9280
rect 3480 9216 3488 9280
rect 3168 8192 3488 9216
rect 3168 8128 3176 8192
rect 3240 8162 3256 8192
rect 3320 8162 3336 8192
rect 3400 8162 3416 8192
rect 3480 8128 3488 8192
rect 3168 7926 3210 8128
rect 3446 7926 3488 8128
rect 3168 7104 3488 7926
rect 3168 7040 3176 7104
rect 3240 7040 3256 7104
rect 3320 7040 3336 7104
rect 3400 7040 3416 7104
rect 3480 7040 3488 7104
rect 3168 6016 3488 7040
rect 3168 5952 3176 6016
rect 3240 5952 3256 6016
rect 3320 5952 3336 6016
rect 3400 5952 3416 6016
rect 3480 5952 3488 6016
rect 3168 4928 3488 5952
rect 3168 4864 3176 4928
rect 3240 4864 3256 4928
rect 3320 4864 3336 4928
rect 3400 4864 3416 4928
rect 3480 4864 3488 4928
rect 3168 4250 3488 4864
rect 3168 4014 3210 4250
rect 3446 4014 3488 4250
rect 3168 3840 3488 4014
rect 3168 3776 3176 3840
rect 3240 3776 3256 3840
rect 3320 3776 3336 3840
rect 3400 3776 3416 3840
rect 3480 3776 3488 3840
rect 3168 2752 3488 3776
rect 3168 2688 3176 2752
rect 3240 2688 3256 2752
rect 3320 2688 3336 2752
rect 3400 2688 3416 2752
rect 3480 2688 3488 2752
rect 3168 2128 3488 2688
rect 5392 17440 5712 17456
rect 5392 17376 5400 17440
rect 5464 17376 5480 17440
rect 5544 17376 5560 17440
rect 5624 17376 5640 17440
rect 5704 17376 5712 17440
rect 5392 16352 5712 17376
rect 5392 16288 5400 16352
rect 5464 16288 5480 16352
rect 5544 16288 5560 16352
rect 5624 16288 5640 16352
rect 5704 16288 5712 16352
rect 5392 15264 5712 16288
rect 5392 15200 5400 15264
rect 5464 15200 5480 15264
rect 5544 15200 5560 15264
rect 5624 15200 5640 15264
rect 5704 15200 5712 15264
rect 5392 14176 5712 15200
rect 5392 14112 5400 14176
rect 5464 14112 5480 14176
rect 5544 14112 5560 14176
rect 5624 14112 5640 14176
rect 5704 14112 5712 14176
rect 5392 14030 5712 14112
rect 5392 13794 5434 14030
rect 5670 13794 5712 14030
rect 5392 13088 5712 13794
rect 5392 13024 5400 13088
rect 5464 13024 5480 13088
rect 5544 13024 5560 13088
rect 5624 13024 5640 13088
rect 5704 13024 5712 13088
rect 5392 12000 5712 13024
rect 5392 11936 5400 12000
rect 5464 11936 5480 12000
rect 5544 11936 5560 12000
rect 5624 11936 5640 12000
rect 5704 11936 5712 12000
rect 5392 10912 5712 11936
rect 5392 10848 5400 10912
rect 5464 10848 5480 10912
rect 5544 10848 5560 10912
rect 5624 10848 5640 10912
rect 5704 10848 5712 10912
rect 5392 10118 5712 10848
rect 5392 9882 5434 10118
rect 5670 9882 5712 10118
rect 5392 9824 5712 9882
rect 5392 9760 5400 9824
rect 5464 9760 5480 9824
rect 5544 9760 5560 9824
rect 5624 9760 5640 9824
rect 5704 9760 5712 9824
rect 5392 8736 5712 9760
rect 5392 8672 5400 8736
rect 5464 8672 5480 8736
rect 5544 8672 5560 8736
rect 5624 8672 5640 8736
rect 5704 8672 5712 8736
rect 5392 7648 5712 8672
rect 5392 7584 5400 7648
rect 5464 7584 5480 7648
rect 5544 7584 5560 7648
rect 5624 7584 5640 7648
rect 5704 7584 5712 7648
rect 5392 6560 5712 7584
rect 5392 6496 5400 6560
rect 5464 6496 5480 6560
rect 5544 6496 5560 6560
rect 5624 6496 5640 6560
rect 5704 6496 5712 6560
rect 5392 6206 5712 6496
rect 5392 5970 5434 6206
rect 5670 5970 5712 6206
rect 5392 5472 5712 5970
rect 5392 5408 5400 5472
rect 5464 5408 5480 5472
rect 5544 5408 5560 5472
rect 5624 5408 5640 5472
rect 5704 5408 5712 5472
rect 5392 4384 5712 5408
rect 5392 4320 5400 4384
rect 5464 4320 5480 4384
rect 5544 4320 5560 4384
rect 5624 4320 5640 4384
rect 5704 4320 5712 4384
rect 5392 3296 5712 4320
rect 5392 3232 5400 3296
rect 5464 3232 5480 3296
rect 5544 3232 5560 3296
rect 5624 3232 5640 3296
rect 5704 3232 5712 3296
rect 5392 2208 5712 3232
rect 5392 2144 5400 2208
rect 5464 2144 5480 2208
rect 5544 2144 5560 2208
rect 5624 2144 5640 2208
rect 5704 2144 5712 2208
rect 5392 2128 5712 2144
rect 7616 16896 7936 17456
rect 7616 16832 7624 16896
rect 7688 16832 7704 16896
rect 7768 16832 7784 16896
rect 7848 16832 7864 16896
rect 7928 16832 7936 16896
rect 7616 15986 7936 16832
rect 7616 15808 7658 15986
rect 7894 15808 7936 15986
rect 7616 15744 7624 15808
rect 7688 15744 7704 15750
rect 7768 15744 7784 15750
rect 7848 15744 7864 15750
rect 7928 15744 7936 15808
rect 7616 14720 7936 15744
rect 7616 14656 7624 14720
rect 7688 14656 7704 14720
rect 7768 14656 7784 14720
rect 7848 14656 7864 14720
rect 7928 14656 7936 14720
rect 7616 13632 7936 14656
rect 7616 13568 7624 13632
rect 7688 13568 7704 13632
rect 7768 13568 7784 13632
rect 7848 13568 7864 13632
rect 7928 13568 7936 13632
rect 7616 12544 7936 13568
rect 7616 12480 7624 12544
rect 7688 12480 7704 12544
rect 7768 12480 7784 12544
rect 7848 12480 7864 12544
rect 7928 12480 7936 12544
rect 7616 12074 7936 12480
rect 7616 11838 7658 12074
rect 7894 11838 7936 12074
rect 7616 11456 7936 11838
rect 7616 11392 7624 11456
rect 7688 11392 7704 11456
rect 7768 11392 7784 11456
rect 7848 11392 7864 11456
rect 7928 11392 7936 11456
rect 7616 10368 7936 11392
rect 7616 10304 7624 10368
rect 7688 10304 7704 10368
rect 7768 10304 7784 10368
rect 7848 10304 7864 10368
rect 7928 10304 7936 10368
rect 7616 9280 7936 10304
rect 7616 9216 7624 9280
rect 7688 9216 7704 9280
rect 7768 9216 7784 9280
rect 7848 9216 7864 9280
rect 7928 9216 7936 9280
rect 7616 8192 7936 9216
rect 7616 8128 7624 8192
rect 7688 8162 7704 8192
rect 7768 8162 7784 8192
rect 7848 8162 7864 8192
rect 7928 8128 7936 8192
rect 7616 7926 7658 8128
rect 7894 7926 7936 8128
rect 7616 7104 7936 7926
rect 7616 7040 7624 7104
rect 7688 7040 7704 7104
rect 7768 7040 7784 7104
rect 7848 7040 7864 7104
rect 7928 7040 7936 7104
rect 7616 6016 7936 7040
rect 7616 5952 7624 6016
rect 7688 5952 7704 6016
rect 7768 5952 7784 6016
rect 7848 5952 7864 6016
rect 7928 5952 7936 6016
rect 7616 4928 7936 5952
rect 7616 4864 7624 4928
rect 7688 4864 7704 4928
rect 7768 4864 7784 4928
rect 7848 4864 7864 4928
rect 7928 4864 7936 4928
rect 7616 4250 7936 4864
rect 7616 4014 7658 4250
rect 7894 4014 7936 4250
rect 7616 3840 7936 4014
rect 7616 3776 7624 3840
rect 7688 3776 7704 3840
rect 7768 3776 7784 3840
rect 7848 3776 7864 3840
rect 7928 3776 7936 3840
rect 7616 2752 7936 3776
rect 7616 2688 7624 2752
rect 7688 2688 7704 2752
rect 7768 2688 7784 2752
rect 7848 2688 7864 2752
rect 7928 2688 7936 2752
rect 7616 2128 7936 2688
rect 9840 17440 10160 17456
rect 9840 17376 9848 17440
rect 9912 17376 9928 17440
rect 9992 17376 10008 17440
rect 10072 17376 10088 17440
rect 10152 17376 10160 17440
rect 9840 16352 10160 17376
rect 9840 16288 9848 16352
rect 9912 16288 9928 16352
rect 9992 16288 10008 16352
rect 10072 16288 10088 16352
rect 10152 16288 10160 16352
rect 9840 15264 10160 16288
rect 9840 15200 9848 15264
rect 9912 15200 9928 15264
rect 9992 15200 10008 15264
rect 10072 15200 10088 15264
rect 10152 15200 10160 15264
rect 9840 14176 10160 15200
rect 9840 14112 9848 14176
rect 9912 14112 9928 14176
rect 9992 14112 10008 14176
rect 10072 14112 10088 14176
rect 10152 14112 10160 14176
rect 9840 14030 10160 14112
rect 9840 13794 9882 14030
rect 10118 13794 10160 14030
rect 9840 13088 10160 13794
rect 9840 13024 9848 13088
rect 9912 13024 9928 13088
rect 9992 13024 10008 13088
rect 10072 13024 10088 13088
rect 10152 13024 10160 13088
rect 9840 12000 10160 13024
rect 9840 11936 9848 12000
rect 9912 11936 9928 12000
rect 9992 11936 10008 12000
rect 10072 11936 10088 12000
rect 10152 11936 10160 12000
rect 9840 10912 10160 11936
rect 9840 10848 9848 10912
rect 9912 10848 9928 10912
rect 9992 10848 10008 10912
rect 10072 10848 10088 10912
rect 10152 10848 10160 10912
rect 9840 10118 10160 10848
rect 9840 9882 9882 10118
rect 10118 9882 10160 10118
rect 9840 9824 10160 9882
rect 9840 9760 9848 9824
rect 9912 9760 9928 9824
rect 9992 9760 10008 9824
rect 10072 9760 10088 9824
rect 10152 9760 10160 9824
rect 9840 8736 10160 9760
rect 9840 8672 9848 8736
rect 9912 8672 9928 8736
rect 9992 8672 10008 8736
rect 10072 8672 10088 8736
rect 10152 8672 10160 8736
rect 9840 7648 10160 8672
rect 9840 7584 9848 7648
rect 9912 7584 9928 7648
rect 9992 7584 10008 7648
rect 10072 7584 10088 7648
rect 10152 7584 10160 7648
rect 9840 6560 10160 7584
rect 9840 6496 9848 6560
rect 9912 6496 9928 6560
rect 9992 6496 10008 6560
rect 10072 6496 10088 6560
rect 10152 6496 10160 6560
rect 9840 6206 10160 6496
rect 9840 5970 9882 6206
rect 10118 5970 10160 6206
rect 9840 5472 10160 5970
rect 9840 5408 9848 5472
rect 9912 5408 9928 5472
rect 9992 5408 10008 5472
rect 10072 5408 10088 5472
rect 10152 5408 10160 5472
rect 9840 4384 10160 5408
rect 9840 4320 9848 4384
rect 9912 4320 9928 4384
rect 9992 4320 10008 4384
rect 10072 4320 10088 4384
rect 10152 4320 10160 4384
rect 9840 3296 10160 4320
rect 9840 3232 9848 3296
rect 9912 3232 9928 3296
rect 9992 3232 10008 3296
rect 10072 3232 10088 3296
rect 10152 3232 10160 3296
rect 9840 2208 10160 3232
rect 9840 2144 9848 2208
rect 9912 2144 9928 2208
rect 9992 2144 10008 2208
rect 10072 2144 10088 2208
rect 10152 2144 10160 2208
rect 9840 2128 10160 2144
rect 12064 16896 12384 17456
rect 12064 16832 12072 16896
rect 12136 16832 12152 16896
rect 12216 16832 12232 16896
rect 12296 16832 12312 16896
rect 12376 16832 12384 16896
rect 12064 15986 12384 16832
rect 12064 15808 12106 15986
rect 12342 15808 12384 15986
rect 12064 15744 12072 15808
rect 12136 15744 12152 15750
rect 12216 15744 12232 15750
rect 12296 15744 12312 15750
rect 12376 15744 12384 15808
rect 12064 14720 12384 15744
rect 12064 14656 12072 14720
rect 12136 14656 12152 14720
rect 12216 14656 12232 14720
rect 12296 14656 12312 14720
rect 12376 14656 12384 14720
rect 12064 13632 12384 14656
rect 12064 13568 12072 13632
rect 12136 13568 12152 13632
rect 12216 13568 12232 13632
rect 12296 13568 12312 13632
rect 12376 13568 12384 13632
rect 12064 12544 12384 13568
rect 12064 12480 12072 12544
rect 12136 12480 12152 12544
rect 12216 12480 12232 12544
rect 12296 12480 12312 12544
rect 12376 12480 12384 12544
rect 12064 12074 12384 12480
rect 12064 11838 12106 12074
rect 12342 11838 12384 12074
rect 12064 11456 12384 11838
rect 12064 11392 12072 11456
rect 12136 11392 12152 11456
rect 12216 11392 12232 11456
rect 12296 11392 12312 11456
rect 12376 11392 12384 11456
rect 12064 10368 12384 11392
rect 12064 10304 12072 10368
rect 12136 10304 12152 10368
rect 12216 10304 12232 10368
rect 12296 10304 12312 10368
rect 12376 10304 12384 10368
rect 12064 9280 12384 10304
rect 12064 9216 12072 9280
rect 12136 9216 12152 9280
rect 12216 9216 12232 9280
rect 12296 9216 12312 9280
rect 12376 9216 12384 9280
rect 12064 8192 12384 9216
rect 12064 8128 12072 8192
rect 12136 8162 12152 8192
rect 12216 8162 12232 8192
rect 12296 8162 12312 8192
rect 12376 8128 12384 8192
rect 12064 7926 12106 8128
rect 12342 7926 12384 8128
rect 12064 7104 12384 7926
rect 12064 7040 12072 7104
rect 12136 7040 12152 7104
rect 12216 7040 12232 7104
rect 12296 7040 12312 7104
rect 12376 7040 12384 7104
rect 12064 6016 12384 7040
rect 12064 5952 12072 6016
rect 12136 5952 12152 6016
rect 12216 5952 12232 6016
rect 12296 5952 12312 6016
rect 12376 5952 12384 6016
rect 12064 4928 12384 5952
rect 12064 4864 12072 4928
rect 12136 4864 12152 4928
rect 12216 4864 12232 4928
rect 12296 4864 12312 4928
rect 12376 4864 12384 4928
rect 12064 4250 12384 4864
rect 12064 4014 12106 4250
rect 12342 4014 12384 4250
rect 12064 3840 12384 4014
rect 12064 3776 12072 3840
rect 12136 3776 12152 3840
rect 12216 3776 12232 3840
rect 12296 3776 12312 3840
rect 12376 3776 12384 3840
rect 12064 2752 12384 3776
rect 12064 2688 12072 2752
rect 12136 2688 12152 2752
rect 12216 2688 12232 2752
rect 12296 2688 12312 2752
rect 12376 2688 12384 2752
rect 12064 2128 12384 2688
rect 14288 17440 14608 17456
rect 14288 17376 14296 17440
rect 14360 17376 14376 17440
rect 14440 17376 14456 17440
rect 14520 17376 14536 17440
rect 14600 17376 14608 17440
rect 14288 16352 14608 17376
rect 14288 16288 14296 16352
rect 14360 16288 14376 16352
rect 14440 16288 14456 16352
rect 14520 16288 14536 16352
rect 14600 16288 14608 16352
rect 14288 15264 14608 16288
rect 14288 15200 14296 15264
rect 14360 15200 14376 15264
rect 14440 15200 14456 15264
rect 14520 15200 14536 15264
rect 14600 15200 14608 15264
rect 14288 14176 14608 15200
rect 14288 14112 14296 14176
rect 14360 14112 14376 14176
rect 14440 14112 14456 14176
rect 14520 14112 14536 14176
rect 14600 14112 14608 14176
rect 14288 14030 14608 14112
rect 14288 13794 14330 14030
rect 14566 13794 14608 14030
rect 14288 13088 14608 13794
rect 14288 13024 14296 13088
rect 14360 13024 14376 13088
rect 14440 13024 14456 13088
rect 14520 13024 14536 13088
rect 14600 13024 14608 13088
rect 14288 12000 14608 13024
rect 14288 11936 14296 12000
rect 14360 11936 14376 12000
rect 14440 11936 14456 12000
rect 14520 11936 14536 12000
rect 14600 11936 14608 12000
rect 14288 10912 14608 11936
rect 14288 10848 14296 10912
rect 14360 10848 14376 10912
rect 14440 10848 14456 10912
rect 14520 10848 14536 10912
rect 14600 10848 14608 10912
rect 14288 10118 14608 10848
rect 14288 9882 14330 10118
rect 14566 9882 14608 10118
rect 14288 9824 14608 9882
rect 14288 9760 14296 9824
rect 14360 9760 14376 9824
rect 14440 9760 14456 9824
rect 14520 9760 14536 9824
rect 14600 9760 14608 9824
rect 14288 8736 14608 9760
rect 14288 8672 14296 8736
rect 14360 8672 14376 8736
rect 14440 8672 14456 8736
rect 14520 8672 14536 8736
rect 14600 8672 14608 8736
rect 14288 7648 14608 8672
rect 14288 7584 14296 7648
rect 14360 7584 14376 7648
rect 14440 7584 14456 7648
rect 14520 7584 14536 7648
rect 14600 7584 14608 7648
rect 14288 6560 14608 7584
rect 14288 6496 14296 6560
rect 14360 6496 14376 6560
rect 14440 6496 14456 6560
rect 14520 6496 14536 6560
rect 14600 6496 14608 6560
rect 14288 6206 14608 6496
rect 14288 5970 14330 6206
rect 14566 5970 14608 6206
rect 14288 5472 14608 5970
rect 14288 5408 14296 5472
rect 14360 5408 14376 5472
rect 14440 5408 14456 5472
rect 14520 5408 14536 5472
rect 14600 5408 14608 5472
rect 14288 4384 14608 5408
rect 14288 4320 14296 4384
rect 14360 4320 14376 4384
rect 14440 4320 14456 4384
rect 14520 4320 14536 4384
rect 14600 4320 14608 4384
rect 14288 3296 14608 4320
rect 14288 3232 14296 3296
rect 14360 3232 14376 3296
rect 14440 3232 14456 3296
rect 14520 3232 14536 3296
rect 14600 3232 14608 3296
rect 14288 2208 14608 3232
rect 14288 2144 14296 2208
rect 14360 2144 14376 2208
rect 14440 2144 14456 2208
rect 14520 2144 14536 2208
rect 14600 2144 14608 2208
rect 14288 2128 14608 2144
rect 16512 16896 16832 17456
rect 16512 16832 16520 16896
rect 16584 16832 16600 16896
rect 16664 16832 16680 16896
rect 16744 16832 16760 16896
rect 16824 16832 16832 16896
rect 16512 15986 16832 16832
rect 16512 15808 16554 15986
rect 16790 15808 16832 15986
rect 16512 15744 16520 15808
rect 16584 15744 16600 15750
rect 16664 15744 16680 15750
rect 16744 15744 16760 15750
rect 16824 15744 16832 15808
rect 16512 14720 16832 15744
rect 16512 14656 16520 14720
rect 16584 14656 16600 14720
rect 16664 14656 16680 14720
rect 16744 14656 16760 14720
rect 16824 14656 16832 14720
rect 16512 13632 16832 14656
rect 16512 13568 16520 13632
rect 16584 13568 16600 13632
rect 16664 13568 16680 13632
rect 16744 13568 16760 13632
rect 16824 13568 16832 13632
rect 16512 12544 16832 13568
rect 16512 12480 16520 12544
rect 16584 12480 16600 12544
rect 16664 12480 16680 12544
rect 16744 12480 16760 12544
rect 16824 12480 16832 12544
rect 16512 12074 16832 12480
rect 16512 11838 16554 12074
rect 16790 11838 16832 12074
rect 16512 11456 16832 11838
rect 16512 11392 16520 11456
rect 16584 11392 16600 11456
rect 16664 11392 16680 11456
rect 16744 11392 16760 11456
rect 16824 11392 16832 11456
rect 16512 10368 16832 11392
rect 16512 10304 16520 10368
rect 16584 10304 16600 10368
rect 16664 10304 16680 10368
rect 16744 10304 16760 10368
rect 16824 10304 16832 10368
rect 16512 9280 16832 10304
rect 16512 9216 16520 9280
rect 16584 9216 16600 9280
rect 16664 9216 16680 9280
rect 16744 9216 16760 9280
rect 16824 9216 16832 9280
rect 16512 8192 16832 9216
rect 16512 8128 16520 8192
rect 16584 8162 16600 8192
rect 16664 8162 16680 8192
rect 16744 8162 16760 8192
rect 16824 8128 16832 8192
rect 16512 7926 16554 8128
rect 16790 7926 16832 8128
rect 16512 7104 16832 7926
rect 16512 7040 16520 7104
rect 16584 7040 16600 7104
rect 16664 7040 16680 7104
rect 16744 7040 16760 7104
rect 16824 7040 16832 7104
rect 16512 6016 16832 7040
rect 16512 5952 16520 6016
rect 16584 5952 16600 6016
rect 16664 5952 16680 6016
rect 16744 5952 16760 6016
rect 16824 5952 16832 6016
rect 16512 4928 16832 5952
rect 16512 4864 16520 4928
rect 16584 4864 16600 4928
rect 16664 4864 16680 4928
rect 16744 4864 16760 4928
rect 16824 4864 16832 4928
rect 16512 4250 16832 4864
rect 16512 4014 16554 4250
rect 16790 4014 16832 4250
rect 16512 3840 16832 4014
rect 16512 3776 16520 3840
rect 16584 3776 16600 3840
rect 16664 3776 16680 3840
rect 16744 3776 16760 3840
rect 16824 3776 16832 3840
rect 16512 2752 16832 3776
rect 16512 2688 16520 2752
rect 16584 2688 16600 2752
rect 16664 2688 16680 2752
rect 16744 2688 16760 2752
rect 16824 2688 16832 2752
rect 16512 2128 16832 2688
<< via4 >>
rect 3210 15808 3446 15986
rect 3210 15750 3240 15808
rect 3240 15750 3256 15808
rect 3256 15750 3320 15808
rect 3320 15750 3336 15808
rect 3336 15750 3400 15808
rect 3400 15750 3416 15808
rect 3416 15750 3446 15808
rect 3210 11838 3446 12074
rect 3210 8128 3240 8162
rect 3240 8128 3256 8162
rect 3256 8128 3320 8162
rect 3320 8128 3336 8162
rect 3336 8128 3400 8162
rect 3400 8128 3416 8162
rect 3416 8128 3446 8162
rect 3210 7926 3446 8128
rect 3210 4014 3446 4250
rect 5434 13794 5670 14030
rect 5434 9882 5670 10118
rect 5434 5970 5670 6206
rect 7658 15808 7894 15986
rect 7658 15750 7688 15808
rect 7688 15750 7704 15808
rect 7704 15750 7768 15808
rect 7768 15750 7784 15808
rect 7784 15750 7848 15808
rect 7848 15750 7864 15808
rect 7864 15750 7894 15808
rect 7658 11838 7894 12074
rect 7658 8128 7688 8162
rect 7688 8128 7704 8162
rect 7704 8128 7768 8162
rect 7768 8128 7784 8162
rect 7784 8128 7848 8162
rect 7848 8128 7864 8162
rect 7864 8128 7894 8162
rect 7658 7926 7894 8128
rect 7658 4014 7894 4250
rect 9882 13794 10118 14030
rect 9882 9882 10118 10118
rect 9882 5970 10118 6206
rect 12106 15808 12342 15986
rect 12106 15750 12136 15808
rect 12136 15750 12152 15808
rect 12152 15750 12216 15808
rect 12216 15750 12232 15808
rect 12232 15750 12296 15808
rect 12296 15750 12312 15808
rect 12312 15750 12342 15808
rect 12106 11838 12342 12074
rect 12106 8128 12136 8162
rect 12136 8128 12152 8162
rect 12152 8128 12216 8162
rect 12216 8128 12232 8162
rect 12232 8128 12296 8162
rect 12296 8128 12312 8162
rect 12312 8128 12342 8162
rect 12106 7926 12342 8128
rect 12106 4014 12342 4250
rect 14330 13794 14566 14030
rect 14330 9882 14566 10118
rect 14330 5970 14566 6206
rect 16554 15808 16790 15986
rect 16554 15750 16584 15808
rect 16584 15750 16600 15808
rect 16600 15750 16664 15808
rect 16664 15750 16680 15808
rect 16680 15750 16744 15808
rect 16744 15750 16760 15808
rect 16760 15750 16790 15808
rect 16554 11838 16790 12074
rect 16554 8128 16584 8162
rect 16584 8128 16600 8162
rect 16600 8128 16664 8162
rect 16664 8128 16680 8162
rect 16680 8128 16744 8162
rect 16744 8128 16760 8162
rect 16760 8128 16790 8162
rect 16554 7926 16790 8128
rect 16554 4014 16790 4250
<< metal5 >>
rect 1056 15986 18908 16028
rect 1056 15750 3210 15986
rect 3446 15750 7658 15986
rect 7894 15750 12106 15986
rect 12342 15750 16554 15986
rect 16790 15750 18908 15986
rect 1056 15708 18908 15750
rect 1056 14030 18908 14072
rect 1056 13794 5434 14030
rect 5670 13794 9882 14030
rect 10118 13794 14330 14030
rect 14566 13794 18908 14030
rect 1056 13752 18908 13794
rect 1056 12074 18908 12116
rect 1056 11838 3210 12074
rect 3446 11838 7658 12074
rect 7894 11838 12106 12074
rect 12342 11838 16554 12074
rect 16790 11838 18908 12074
rect 1056 11796 18908 11838
rect 1056 10118 18908 10160
rect 1056 9882 5434 10118
rect 5670 9882 9882 10118
rect 10118 9882 14330 10118
rect 14566 9882 18908 10118
rect 1056 9840 18908 9882
rect 1056 8162 18908 8204
rect 1056 7926 3210 8162
rect 3446 7926 7658 8162
rect 7894 7926 12106 8162
rect 12342 7926 16554 8162
rect 16790 7926 18908 8162
rect 1056 7884 18908 7926
rect 1056 6206 18908 6248
rect 1056 5970 5434 6206
rect 5670 5970 9882 6206
rect 10118 5970 14330 6206
rect 14566 5970 18908 6206
rect 1056 5928 18908 5970
rect 1056 4250 18908 4292
rect 1056 4014 3210 4250
rect 3446 4014 7658 4250
rect 7894 4014 12106 4250
rect 12342 4014 16554 4250
rect 16790 4014 18908 4250
rect 1056 3972 18908 4014
use sky130_ef_sc_hd__decap_12  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1649977179
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1649977179
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1649977179
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1649977179
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1649977179
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1649977179
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1649977179
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1649977179
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1649977179
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1649977179
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1649977179
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1649977179
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1649977179
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_153 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 15180 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_161 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 15916 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_167
timestamp 1649977179
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1649977179
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_181 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 17756 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_189
timestamp 1649977179
transform 1 0 18492 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1649977179
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1649977179
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1649977179
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1649977179
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1649977179
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1649977179
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1649977179
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1649977179
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1649977179
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1649977179
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1649977179
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1649977179
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1649977179
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1649977179
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1649977179
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1649977179
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1649977179
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1649977179
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1649977179
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_181
timestamp 1649977179
transform 1 0 17756 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_189
timestamp 1649977179
transform 1 0 18492 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1649977179
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1649977179
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1649977179
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1649977179
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1649977179
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1649977179
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1649977179
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1649977179
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1649977179
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1649977179
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1649977179
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1649977179
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1649977179
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1649977179
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1649977179
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1649977179
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1649977179
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1649977179
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1649977179
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_189
timestamp 1649977179
transform 1 0 18492 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1649977179
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1649977179
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1649977179
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1649977179
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1649977179
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1649977179
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1649977179
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1649977179
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1649977179
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1649977179
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1649977179
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1649977179
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1649977179
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1649977179
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1649977179
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1649977179
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1649977179
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1649977179
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1649977179
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_181
timestamp 1649977179
transform 1 0 17756 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_189
timestamp 1649977179
transform 1 0 18492 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1649977179
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1649977179
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1649977179
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1649977179
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1649977179
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1649977179
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1649977179
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1649977179
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1649977179
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1649977179
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1649977179
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1649977179
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1649977179
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1649977179
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1649977179
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1649977179
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1649977179
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1649977179
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1649977179
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_189
timestamp 1649977179
transform 1 0 18492 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1649977179
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1649977179
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1649977179
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1649977179
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1649977179
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1649977179
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1649977179
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1649977179
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1649977179
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1649977179
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1649977179
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1649977179
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1649977179
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1649977179
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1649977179
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1649977179
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1649977179
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1649977179
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1649977179
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_181
timestamp 1649977179
transform 1 0 17756 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_189
timestamp 1649977179
transform 1 0 18492 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1649977179
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1649977179
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1649977179
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1649977179
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1649977179
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1649977179
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1649977179
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1649977179
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1649977179
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1649977179
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1649977179
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1649977179
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1649977179
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1649977179
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1649977179
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1649977179
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1649977179
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1649977179
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1649977179
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_189
timestamp 1649977179
transform 1 0 18492 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1649977179
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1649977179
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1649977179
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1649977179
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1649977179
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1649977179
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1649977179
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1649977179
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1649977179
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1649977179
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1649977179
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1649977179
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1649977179
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1649977179
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1649977179
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1649977179
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1649977179
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1649977179
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1649977179
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_181
timestamp 1649977179
transform 1 0 17756 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_189
timestamp 1649977179
transform 1 0 18492 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1649977179
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1649977179
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1649977179
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1649977179
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1649977179
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1649977179
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1649977179
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1649977179
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1649977179
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1649977179
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1649977179
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1649977179
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1649977179
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1649977179
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1649977179
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1649977179
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1649977179
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1649977179
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1649977179
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_189
timestamp 1649977179
transform 1 0 18492 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1649977179
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1649977179
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1649977179
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1649977179
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1649977179
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1649977179
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1649977179
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1649977179
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1649977179
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1649977179
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1649977179
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1649977179
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1649977179
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1649977179
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1649977179
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1649977179
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1649977179
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1649977179
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1649977179
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_181
timestamp 1649977179
transform 1 0 17756 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_189
timestamp 1649977179
transform 1 0 18492 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1649977179
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1649977179
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1649977179
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1649977179
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1649977179
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1649977179
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1649977179
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1649977179
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1649977179
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1649977179
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_97
timestamp 1649977179
transform 1 0 10028 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1649977179
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1649977179
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1649977179
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1649977179
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1649977179
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1649977179
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1649977179
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_189
timestamp 1649977179
transform 1 0 18492 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1649977179
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1649977179
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1649977179
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1649977179
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1649977179
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1649977179
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1649977179
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1649977179
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1649977179
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1649977179
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1649977179
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1649977179
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1649977179
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1649977179
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1649977179
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1649977179
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1649977179
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1649977179
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1649977179
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_181
timestamp 1649977179
transform 1 0 17756 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_189
timestamp 1649977179
transform 1 0 18492 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1649977179
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1649977179
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1649977179
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1649977179
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1649977179
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1649977179
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1649977179
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1649977179
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1649977179
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1649977179
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1649977179
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1649977179
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1649977179
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1649977179
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1649977179
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1649977179
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1649977179
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1649977179
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1649977179
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_189
timestamp 1649977179
transform 1 0 18492 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1649977179
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1649977179
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1649977179
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1649977179
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1649977179
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1649977179
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1649977179
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1649977179
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1649977179
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1649977179
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1649977179
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1649977179
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1649977179
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1649977179
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1649977179
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1649977179
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1649977179
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1649977179
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1649977179
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_181
timestamp 1649977179
transform 1 0 17756 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_189
timestamp 1649977179
transform 1 0 18492 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1649977179
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1649977179
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1649977179
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1649977179
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1649977179
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1649977179
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1649977179
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1649977179
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1649977179
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1649977179
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1649977179
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_109
timestamp 1649977179
transform 1 0 11132 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_129
timestamp 1649977179
transform 1 0 12972 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_137
timestamp 1649977179
transform 1 0 13708 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1649977179
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1649977179
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_165
timestamp 1649977179
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_177
timestamp 1649977179
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_189
timestamp 1649977179
transform 1 0 18492 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1649977179
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1649977179
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1649977179
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1649977179
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1649977179
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1649977179
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1649977179
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_69
timestamp 1649977179
transform 1 0 7452 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1649977179
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1649977179
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1649977179
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_129
timestamp 1649977179
transform 1 0 12972 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_141
timestamp 1649977179
transform 1 0 14076 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_153
timestamp 1649977179
transform 1 0 15180 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_165
timestamp 1649977179
transform 1 0 16284 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1649977179
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_181
timestamp 1649977179
transform 1 0 17756 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_189
timestamp 1649977179
transform 1 0 18492 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1649977179
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1649977179
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1649977179
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1649977179
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1649977179
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1649977179
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1649977179
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1649977179
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1649977179
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1649977179
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1649977179
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_109
timestamp 1649977179
transform 1 0 11132 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_132
timestamp 1649977179
transform 1 0 13248 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_16_147
timestamp 1649977179
transform 1 0 14628 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_159
timestamp 1649977179
transform 1 0 15732 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_171
timestamp 1649977179
transform 1 0 16836 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_183
timestamp 1649977179
transform 1 0 17940 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_189
timestamp 1649977179
transform 1 0 18492 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1649977179
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1649977179
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1649977179
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1649977179
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1649977179
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1649977179
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1649977179
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1649977179
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1649977179
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_93
timestamp 1649977179
transform 1 0 9660 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_108
timestamp 1649977179
transform 1 0 11040 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_121
timestamp 1649977179
transform 1 0 12236 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_128
timestamp 1649977179
transform 1 0 12880 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_140
timestamp 1649977179
transform 1 0 13984 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_152
timestamp 1649977179
transform 1 0 15088 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_164
timestamp 1649977179
transform 1 0 16192 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1649977179
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_181 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 17756 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_186
timestamp 1649977179
transform 1 0 18216 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1649977179
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1649977179
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1649977179
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1649977179
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1649977179
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1649977179
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1649977179
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1649977179
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1649977179
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1649977179
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1649977179
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_109
timestamp 1649977179
transform 1 0 11132 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_119
timestamp 1649977179
transform 1 0 12052 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_131
timestamp 1649977179
transform 1 0 13156 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1649977179
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1649977179
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_153
timestamp 1649977179
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_165
timestamp 1649977179
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_177
timestamp 1649977179
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_189
timestamp 1649977179
transform 1 0 18492 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1649977179
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1649977179
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1649977179
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1649977179
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1649977179
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1649977179
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1649977179
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1649977179
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1649977179
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1649977179
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1649977179
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1649977179
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1649977179
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1649977179
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_137
timestamp 1649977179
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_149
timestamp 1649977179
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1649977179
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1649977179
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1649977179
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_181
timestamp 1649977179
transform 1 0 17756 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_189
timestamp 1649977179
transform 1 0 18492 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1649977179
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1649977179
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1649977179
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1649977179
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1649977179
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1649977179
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1649977179
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1649977179
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1649977179
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1649977179
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1649977179
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1649977179
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_121
timestamp 1649977179
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1649977179
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1649977179
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1649977179
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_153
timestamp 1649977179
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_165
timestamp 1649977179
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_177
timestamp 1649977179
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_189
timestamp 1649977179
transform 1 0 18492 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1649977179
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1649977179
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1649977179
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 1649977179
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1649977179
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1649977179
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1649977179
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1649977179
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1649977179
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1649977179
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1649977179
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1649977179
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1649977179
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_125
timestamp 1649977179
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_137
timestamp 1649977179
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_149
timestamp 1649977179
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1649977179
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1649977179
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1649977179
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_181
timestamp 1649977179
transform 1 0 17756 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_189
timestamp 1649977179
transform 1 0 18492 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1649977179
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1649977179
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1649977179
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1649977179
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1649977179
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1649977179
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1649977179
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1649977179
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1649977179
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1649977179
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1649977179
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_109
timestamp 1649977179
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_121
timestamp 1649977179
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1649977179
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1649977179
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1649977179
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_153
timestamp 1649977179
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_165
timestamp 1649977179
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_177
timestamp 1649977179
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_189
timestamp 1649977179
transform 1 0 18492 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1649977179
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1649977179
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1649977179
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1649977179
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1649977179
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1649977179
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1649977179
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1649977179
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1649977179
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1649977179
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1649977179
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1649977179
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1649977179
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1649977179
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 1649977179
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_149
timestamp 1649977179
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1649977179
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1649977179
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1649977179
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_181
timestamp 1649977179
transform 1 0 17756 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_189
timestamp 1649977179
transform 1 0 18492 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1649977179
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1649977179
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1649977179
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1649977179
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1649977179
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1649977179
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1649977179
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1649977179
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1649977179
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1649977179
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1649977179
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1649977179
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 1649977179
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1649977179
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1649977179
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1649977179
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_153
timestamp 1649977179
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_165
timestamp 1649977179
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_177
timestamp 1649977179
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_189
timestamp 1649977179
transform 1 0 18492 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1649977179
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1649977179
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1649977179
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_39
timestamp 1649977179
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1649977179
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1649977179
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1649977179
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1649977179
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1649977179
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 1649977179
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1649977179
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1649977179
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1649977179
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1649977179
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_137
timestamp 1649977179
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_149
timestamp 1649977179
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1649977179
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1649977179
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1649977179
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_181
timestamp 1649977179
transform 1 0 17756 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_189
timestamp 1649977179
transform 1 0 18492 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_6
timestamp 1649977179
transform 1 0 1656 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_18
timestamp 1649977179
transform 1 0 2760 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_26
timestamp 1649977179
transform 1 0 3496 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1649977179
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1649977179
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1649977179
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1649977179
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1649977179
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1649977179
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1649977179
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1649977179
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1649977179
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_121
timestamp 1649977179
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1649977179
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1649977179
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1649977179
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1649977179
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_165
timestamp 1649977179
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_177
timestamp 1649977179
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_189
timestamp 1649977179
transform 1 0 18492 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1649977179
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1649977179
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_27
timestamp 1649977179
transform 1 0 3588 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_29
timestamp 1649977179
transform 1 0 3772 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_41
timestamp 1649977179
transform 1 0 4876 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_53
timestamp 1649977179
transform 1 0 5980 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1649977179
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1649977179
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_81
timestamp 1649977179
transform 1 0 8556 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_85
timestamp 1649977179
transform 1 0 8924 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_97
timestamp 1649977179
transform 1 0 10028 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_109
timestamp 1649977179
transform 1 0 11132 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_113
timestamp 1649977179
transform 1 0 11500 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_118
timestamp 1649977179
transform 1 0 11960 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_130
timestamp 1649977179
transform 1 0 13064 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_138
timestamp 1649977179
transform 1 0 13800 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_141
timestamp 1649977179
transform 1 0 14076 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_153
timestamp 1649977179
transform 1 0 15180 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_165
timestamp 1649977179
transform 1 0 16284 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 1649977179
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_181
timestamp 1649977179
transform 1 0 17756 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_189
timestamp 1649977179
transform 1 0 18492 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 18860 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 18860 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 18860 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 18860 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 18860 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 18860 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 18860 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 18860 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 18860 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 18860 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 18860 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 18860 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 18860 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 18860 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 18860 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 18860 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 18860 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 18860 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 18860 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 18860 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 18860 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1649977179
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1649977179
transform -1 0 18860 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1649977179
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1649977179
transform -1 0 18860 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1649977179
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1649977179
transform -1 0 18860 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1649977179
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1649977179
transform -1 0 18860 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1649977179
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1649977179
transform -1 0 18860 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1649977179
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1649977179
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1649977179
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1649977179
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1649977179
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1649977179
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1649977179
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1649977179
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1649977179
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1649977179
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1649977179
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1649977179
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1649977179
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1649977179
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1649977179
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1649977179
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1649977179
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1649977179
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1649977179
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1649977179
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1649977179
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1649977179
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1649977179
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1649977179
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1649977179
transform 1 0 3680 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1649977179
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1649977179
transform 1 0 8832 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1649977179
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1649977179
transform 1 0 13984 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1649977179
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _05_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 12880 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _06_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 10396 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _07_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 11316 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__and4b_1  _08_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 11500 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _09_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 14076 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _10_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 11500 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _11_
timestamp 1649977179
transform 1 0 11500 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 11408 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1649977179
transform 1 0 10396 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1649977179
transform -1 0 9660 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 1656 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1649977179
transform 1 0 17940 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1649977179
transform -1 0 11960 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output4 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 15548 0 1 2176
box -38 -48 406 592
<< labels >>
flabel metal4 s 5392 2128 5712 17456 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 9840 2128 10160 17456 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 14288 2128 14608 17456 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 5928 18908 6248 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 9840 18908 10160 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 13752 18908 14072 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 3168 2128 3488 17456 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 7616 2128 7936 17456 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 12064 2128 12384 17456 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 16512 2128 16832 17456 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 3972 18908 4292 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 7884 18908 8204 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 11796 18908 12116 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 15708 18908 16028 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 16328 800 16448 0 FreeSans 480 0 0 0 a
port 2 nsew signal input
flabel metal2 s 18 0 74 800 0 FreeSans 224 90 0 0 clk
port 3 nsew signal input
flabel metal3 s 19200 11568 20000 11688 0 FreeSans 480 0 0 0 en
port 4 nsew signal input
flabel metal2 s 11610 19200 11666 20000 0 FreeSans 224 90 0 0 reset
port 5 nsew signal input
flabel metal2 s 15474 0 15530 800 0 FreeSans 224 90 0 0 y
port 6 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 20000 20000
<< end >>
