module tm1638_led_display_keys
(
    input   clk,
    input   rst,
    output  out_clk,
    output  out_stb,
    input   iodata
);

endmodule
